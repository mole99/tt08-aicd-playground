** sch_path: /home/leo/Projects/tt08-aicd-playground/xschem/tt_um_tt08_aicd_playground.sch
.subckt tt_um_tt08_aicd_playground VAPWR ui_in[7] ui_in[6] ui_in[5] ui_in[4] ui_in[3] ui_in[2] ui_in[1] ui_in[0] VDPWR VGND
+ uio_in[7] uio_in[6] uio_in[5] uio_in[4] uio_in[3] uio_in[2] uio_in[1] uio_in[0] ena uo_out[7] uo_out[6] uo_out[5] uo_out[4] uo_out[3]
+ uo_out[2] uo_out[1] uo_out[0] clk rst_n uio_out[7] uio_out[6] uio_out[5] uio_out[4] uio_out[3] uio_out[2] uio_out[1] uio_out[0] uio_oe[7]
+ uio_oe[6] uio_oe[5] uio_oe[4] uio_oe[3] uio_oe[2] uio_oe[1] uio_oe[0] ua[7] ua[6] ua[5] ua[4] ua[3] ua[2] ua[1] ua[0]
*.PININFO ui_in[7:0]:I uo_out[7:0]:O VGND:B VDPWR:B VAPWR:B uio_in[7:0]:I ua[7:0]:B uio_out[7:0]:O uio_oe[7:0]:O ena:I clk:I
*+ rst_n:I
x1 VDPWR VGND clk net2 ena port_ms_i port_ms_o[0] port_ms_o[1] port_ms_o[2] port_ms_o[3] port_ms_o[4] port_ms_o[5] port_ms_o[6]
+ port_ms_o[7] rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4]
+ uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1]
+ uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6] uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6]
+ uo_out[7] dig_ctrl_top
* noconn ua[7:2]
* noconn #net3
x2[7] VAPWR VDPWR port_ms_o_ana[7] port_ms_o[7] VGND sky130_leo_ip__levelshifter_up
x2[6] VAPWR VDPWR port_ms_o_ana[6] port_ms_o[6] VGND sky130_leo_ip__levelshifter_up
x2[5] VAPWR VDPWR port_ms_o_ana[5] port_ms_o[5] VGND sky130_leo_ip__levelshifter_up
x2[4] VAPWR VDPWR port_ms_o_ana[4] port_ms_o[4] VGND sky130_leo_ip__levelshifter_up
x2[3] VAPWR VDPWR port_ms_o_ana[3] port_ms_o[3] VGND sky130_leo_ip__levelshifter_up
x2[2] VAPWR VDPWR port_ms_o_ana[2] port_ms_o[2] VGND sky130_leo_ip__levelshifter_up
x2[1] VAPWR VDPWR port_ms_o_ana[1] port_ms_o[1] VGND sky130_leo_ip__levelshifter_up
x2[0] VAPWR VDPWR port_ms_o_ana[0] port_ms_o[0] VGND sky130_leo_ip__levelshifter_up
x3 VDPWR port_ms_i net1 VGND sky130_leo_ip__levelshifter_down
x2 D[0] ua[1] D[1] D[2] D[3] D[4] D[5] D[6] D[7] VGND sky130_leo_ip__rdac_8bit
x1[7] port_ms_o_ana[7] VGND VGND VAPWR VAPWR D[7] sky130_fd_sc_hvl__buf_4
x1[6] port_ms_o_ana[6] VGND VGND VAPWR VAPWR D[6] sky130_fd_sc_hvl__buf_4
x1[5] port_ms_o_ana[5] VGND VGND VAPWR VAPWR D[5] sky130_fd_sc_hvl__buf_4
x1[4] port_ms_o_ana[4] VGND VGND VAPWR VAPWR D[4] sky130_fd_sc_hvl__buf_4
x1[3] port_ms_o_ana[3] VGND VGND VAPWR VAPWR D[3] sky130_fd_sc_hvl__buf_4
x1[2] port_ms_o_ana[2] VGND VGND VAPWR VAPWR D[2] sky130_fd_sc_hvl__buf_4
x1[1] port_ms_o_ana[1] VGND VGND VAPWR VAPWR D[1] sky130_fd_sc_hvl__buf_4
x1[0] port_ms_o_ana[0] VGND VGND VAPWR VAPWR D[0] sky130_fd_sc_hvl__buf_4
x4 VAPWR ua[0] net1 ua[1] VGND net2 net3 sky130_leo_ip__comparator
.ends

* expanding   symbol:  dig_ctrl_top.sym # of pins=13
** sym_path: /home/leo/Projects/tt08-aicd-playground/dependencies/dig_ctrl/xschem/dig_ctrl_top.sym
.include /home/leo/Projects/tt08-aicd-playground/dependencies/dig_ctrl/xschem/../spice/dig_ctrl_top.spice

* expanding   symbol:  sky130_leo_ip__levelshifter_up.sym # of pins=5
** sym_path: /home/leo/Projects/tt08-aicd-playground/dependencies/sky130_leo_ip__levelshifter/xschem/sky130_leo_ip__levelshifter_up.sym
** sch_path: /home/leo/Projects/tt08-aicd-playground/dependencies/sky130_leo_ip__levelshifter/xschem/sky130_leo_ip__levelshifter_up.sch
.subckt sky130_leo_ip__levelshifter_up VDDOUT VDDIN OUT IN VGND
*.PININFO IN:I VGND:B VDDIN:B OUT:O VDDOUT:B
XM1 ctrl_n IN VGND VGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 ctrl_n IN VDDIN VDDIN sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 ctrl ctrl_n VGND VGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 ctrl ctrl_n VDDIN VDDIN sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 OUT p1 VDDOUT VDDOUT sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 p1 ctrl VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM7 p1 OUT VDDOUT VDDOUT sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM8 OUT ctrl_n VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  sky130_leo_ip__levelshifter_down.sym # of pins=4
** sym_path: /home/leo/Projects/tt08-aicd-playground/dependencies/sky130_leo_ip__levelshifter/xschem/sky130_leo_ip__levelshifter_down.sym
** sch_path: /home/leo/Projects/tt08-aicd-playground/dependencies/sky130_leo_ip__levelshifter/xschem/sky130_leo_ip__levelshifter_down.sch
.subckt sky130_leo_ip__levelshifter_down VDDOUT OUT IN VGND
*.PININFO IN:I VGND:B OUT:O VDDOUT:B
XM3 OUT n VGND VGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 OUT n VDDOUT VDDOUT sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 n IN VDDOUT VDDOUT sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 n IN VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  sky130_leo_ip__rdac_8bit.sym # of pins=10
** sym_path: /home/leo/Projects/tt08-aicd-playground/dependencies/sky130_leo_ip__rdac_8bit/xschem/sky130_leo_ip__rdac_8bit.sym
** sch_path: /home/leo/Projects/tt08-aicd-playground/dependencies/sky130_leo_ip__rdac_8bit/xschem/sky130_leo_ip__rdac_8bit.sch
.subckt sky130_leo_ip__rdac_8bit D0 OUT D1 D2 D3 D4 D5 D6 D7 VGND
*.PININFO VGND:B D7:I D6:I D5:I D4:I D3:I D2:I D1:I D0:I OUT:O
**** begin user architecture code


* https://skywater-pdk.readthedocs.io/en/main/rules/device-details.html#p-poly-precision-resistors


**** end user architecture code
XR1 D7 net1 VGND sky130_fd_pr__res_high_po_1p41 L=50 mult=1 m=1
XR2 net1 OUT VGND sky130_fd_pr__res_high_po_1p41 L=50 mult=1 m=1
XR3 OUT net2 VGND sky130_fd_pr__res_high_po_1p41 L=50 mult=1 m=1
XR4 D6 net3 VGND sky130_fd_pr__res_high_po_1p41 L=50 mult=1 m=1
XR5 net3 net2 VGND sky130_fd_pr__res_high_po_1p41 L=50 mult=1 m=1
XR6 net2 net4 VGND sky130_fd_pr__res_high_po_1p41 L=50 mult=1 m=1
XR7 D5 net5 VGND sky130_fd_pr__res_high_po_1p41 L=50 mult=1 m=1
XR8 net5 net4 VGND sky130_fd_pr__res_high_po_1p41 L=50 mult=1 m=1
XR9 net4 net6 VGND sky130_fd_pr__res_high_po_1p41 L=50 mult=1 m=1
XR10 D4 net7 VGND sky130_fd_pr__res_high_po_1p41 L=50 mult=1 m=1
XR11 net7 net6 VGND sky130_fd_pr__res_high_po_1p41 L=50 mult=1 m=1
XR12 net6 net8 VGND sky130_fd_pr__res_high_po_1p41 L=50 mult=1 m=1
XR13 D3 net9 VGND sky130_fd_pr__res_high_po_1p41 L=50 mult=1 m=1
XR14 net9 net8 VGND sky130_fd_pr__res_high_po_1p41 L=50 mult=1 m=1
XR15 net8 net10 VGND sky130_fd_pr__res_high_po_1p41 L=50 mult=1 m=1
XR16 D2 net11 VGND sky130_fd_pr__res_high_po_1p41 L=50 mult=1 m=1
XR17 net11 net10 VGND sky130_fd_pr__res_high_po_1p41 L=50 mult=1 m=1
XR18 net10 net12 VGND sky130_fd_pr__res_high_po_1p41 L=50 mult=1 m=1
XR19 D1 net13 VGND sky130_fd_pr__res_high_po_1p41 L=50 mult=1 m=1
XR20 net13 net12 VGND sky130_fd_pr__res_high_po_1p41 L=50 mult=1 m=1
XR21 net12 net14 VGND sky130_fd_pr__res_high_po_1p41 L=50 mult=1 m=1
XR22 D0 net15 VGND sky130_fd_pr__res_high_po_1p41 L=50 mult=1 m=1
XR23 net15 net14 VGND sky130_fd_pr__res_high_po_1p41 L=50 mult=1 m=1
XR24 net14 net16 VGND sky130_fd_pr__res_high_po_1p41 L=50 mult=1 m=1
XR25 net16 VGND VGND sky130_fd_pr__res_high_po_1p41 L=50 mult=1 m=1
XR26 VGND VGND VGND sky130_fd_pr__res_high_po_1p41 L=50 mult=1 m=1
XR27 VGND VGND VGND sky130_fd_pr__res_high_po_1p41 L=50 mult=1 m=1
.ends


* expanding   symbol:  sky130_leo_ip__comparator.sym # of pins=7
** sym_path: /home/leo/Projects/tt08-aicd-playground/dependencies/sky130_leo_ip__comparator/xschem/sky130_leo_ip__comparator.sym
** sch_path: /home/leo/Projects/tt08-aicd-playground/dependencies/sky130_leo_ip__comparator/xschem/sky130_leo_ip__comparator.sch
.subckt sky130_leo_ip__comparator vdd in_p out_p in_n vss clk out_n
*.PININFO out_n:O in_p:I in_n:I vdd:B vss:B clk:I out_p:O
XR1 vss net2 vss sky130_fd_pr__res_xhigh_po_2p85 L=25 mult=1 m=1
XM7 comp_p comp_n vss vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 net2 net2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 L=5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 comp_n comp_p vss vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 net1 net2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 L=5 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 comp_p in_n net1 vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 comp_n in_p net1 vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 comp_n clk comp_p vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
x1 SR_set_n net4 VSS VSS VDD VDD net3 sky130_fd_sc_hvl__nand2_1
x2 net3 SR_reset_n VSS VSS VDD VDD net4 sky130_fd_sc_hvl__nand2_1
XM8 SR_set_n comp_p vdd vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM9 SR_set_n comp_p vss vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM10 SR_reset_n comp_n vdd vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM11 SR_reset_n comp_n vss vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
x3 net3 VSS VSS VDD VDD out_p sky130_fd_sc_hvl__buf_4
x4 net4 VSS VSS VDD VDD out_n sky130_fd_sc_hvl__buf_4
.ends

.end
