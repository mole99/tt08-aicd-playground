* NGSPICE file created from tt_um_tt08_aicd_playground.ext - technology: sky130A

.subckt sky130_leo_ip__levelshifter_up VDDOUT VDDIN OUT IN VGND
X0 VDDIN a_373_442# a_897_442# VDDIN sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.6 as=0.3 ps=2.6 w=1 l=0.15
X1 OUT a_373_442# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.3 pd=2.6 as=0.3 ps=2.6 w=1 l=0.5
X2 VDDIN IN a_373_442# VDDIN sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.6 as=0.3 ps=2.6 w=1 l=0.15
X3 a_897_442# a_373_442# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.126 ps=1.44 w=0.42 l=0.15
X4 VDDOUT OUT a_1778_346# VDDOUT sky130_fd_pr__pfet_g5v0d10v5 ad=0.126 pd=1.44 as=0.126 ps=1.44 w=0.42 l=0.5
X5 a_1778_346# a_897_442# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.3 pd=2.6 as=0.3 ps=2.6 w=1 l=0.5
X6 VDDOUT a_1778_346# OUT VDDOUT sky130_fd_pr__pfet_g5v0d10v5 ad=0.126 pd=1.44 as=0.126 ps=1.44 w=0.42 l=0.5
X7 a_373_442# IN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.126 ps=1.44 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hvl__buf_4 VGND VNB VPWR VPB X A
X0 a_149_81# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.21 ps=1.78 w=1.5 l=0.5
X1 VGND a_149_81# X VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X2 X a_149_81# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.21375 ps=2.07 w=0.75 l=0.5
X3 X a_149_81# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X4 VPWR a_149_81# X VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X5 a_149_81# A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.105 ps=1.03 w=0.75 l=0.5
X6 VPWR a_149_81# X VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X7 X a_149_81# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.4275 ps=3.57 w=1.5 l=0.5
X8 X a_149_81# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X9 VGND a_149_81# X VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
.ends

.subckt nfet$3 a_60_n40# a_160_0# a_0_0# a_n149_n154#
X0 a_160_0# a_60_n40# a_0_0# a_n149_n154# sky130_fd_pr__nfet_g5v0d10v5 ad=0.3 pd=2.6 as=0.3 ps=2.6 w=1 l=0.5
.ends

.subckt nfet a_90_0# a_48_124# a_n123_n128# a_0_0#
X0 a_90_0# a_48_124# a_0_0# a_n123_n128# sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.126 ps=1.44 w=0.42 l=0.15
.ends

.subckt pfet$3 a_90_0# w_n184_n189# a_0_0# a_48_240#
X0 a_90_0# a_48_240# a_0_0# w_n184_n189# sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.6 as=0.3 ps=2.6 w=1 l=0.15
.ends

.subckt pfet$1 a_60_n40# w_n242_n247# a_160_0# a_0_0#
X0 a_160_0# a_60_n40# a_0_0# w_n242_n247# sky130_fd_pr__pfet_g5v0d10v5 ad=0.126 pd=1.44 as=0.126 ps=1.44 w=0.42 l=0.5
.ends

.subckt sky130_leo_ip__levelshifter_down VDDOUT OUT IN VGND
Xnfet$3_0 IN m1_306_395# VGND VGND nfet$3
Xnfet_0 OUT m1_306_395# VGND VGND nfet
Xpfet$3_0 VDDOUT VDDOUT OUT m1_306_395# pfet$3
Xpfet$1_0 IN VDDOUT VDDOUT m1_306_395# pfet$1
.ends

.subckt sky130_fd_sc_hd__and2_2 VPWR VGND VPB VNB A B X
X0 X a_61_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.16655 ps=1.39 w=1 l=0.15
X1 VPWR a_61_75# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.38 pd=2.76 as=0.195 ps=1.39 w=1 l=0.15
X2 VPWR B a_61_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 VGND B a_147_75# VNB sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 X a_61_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.1118 ps=1.04 w=0.65 l=0.15
X5 VGND a_61_75# X VNB sky130_fd_pr__nfet_01v8 ad=0.247 pd=2.06 as=0.12675 ps=1.04 w=0.65 l=0.15
X6 a_61_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X7 a_147_75# A a_61_75# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__dlclkp_1 VGND VPWR VPB VNB GCLK GATE CLK
X0 a_381_369# GATE VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.09575 pd=0.965 as=0.1664 ps=1.8 w=0.64 l=0.15
X1 a_476_413# a_193_47# a_381_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.09575 ps=0.965 w=0.42 l=0.15
X2 a_957_369# a_642_307# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2032 pd=1.275 as=0.149 ps=1.325 w=0.64 l=0.15
X3 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4 a_1042_47# a_642_307# a_957_369# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 GCLK a_957_369# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.325 w=1 l=0.15
X6 VGND CLK a_1042_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0441 ps=0.63 w=0.42 l=0.15
X7 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 a_651_47# a_193_47# a_476_413# VNB sky130_fd_pr__special_nfet_01v8 ad=0.067125 pd=0.745 as=0.1192 ps=1.09 w=0.39 l=0.15
X9 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10 GCLK a_957_369# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X11 VPWR a_642_307# a_600_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X12 a_476_413# a_27_47# a_396_119# VNB sky130_fd_pr__nfet_01v8 ad=0.1192 pd=1.09 as=0.117125 ps=1.085 w=0.42 l=0.15
X13 VPWR CLK a_957_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.2032 ps=1.275 w=0.64 l=0.15
X14 a_642_307# a_476_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.118125 ps=1.04 w=0.65 l=0.15
X15 a_600_413# a_27_47# a_476_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0987 ps=0.89 w=0.42 l=0.15
X16 VPWR a_476_413# a_642_307# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.27 ps=2.54 w=1 l=0.15
X17 VGND a_642_307# a_651_47# VNB sky130_fd_pr__nfet_01v8 ad=0.118125 pd=1.04 as=0.067125 ps=0.745 w=0.42 l=0.15
X18 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X19 a_396_119# GATE VGND VNB sky130_fd_pr__nfet_01v8 ad=0.117125 pd=1.085 as=0.1281 ps=1.45 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4_2 VPWR VGND VPB VNB B D C A X
X0 a_27_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_27_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_277_297# B a_205_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VPWR A a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.101875 ps=0.99 w=0.65 l=0.15
X5 a_205_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 VPWR a_27_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND a_27_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.19825 pd=1.91 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14825 ps=1.34 w=1 l=0.15
X9 VGND C a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_109_297# D a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X11 VGND A a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__dlxtp_1 VGND VPWR VPB VNB Q D GATE
X0 VPWR D a_299_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1 a_560_47# a_193_47# a_465_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.066 ps=0.745 w=0.36 l=0.15
X2 VGND a_713_21# a_659_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0936 pd=1.24 as=0.0486 ps=0.63 w=0.36 l=0.15
X3 Q a_713_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.092625 ps=0.935 w=0.65 l=0.15
X4 a_465_47# a_299_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X5 VPWR GATE a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X6 a_659_47# a_27_47# a_560_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0486 pd=0.63 as=0.0621 ps=0.705 w=0.36 l=0.15
X7 VGND a_560_47# a_713_21# VNB sky130_fd_pr__nfet_01v8 ad=0.092625 pd=0.935 as=0.169 ps=1.82 w=0.65 l=0.15
X8 VPWR a_713_21# a_644_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.07245 ps=0.765 w=0.42 l=0.15
X9 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 VPWR a_560_47# a_713_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1425 pd=1.285 as=0.26 ps=2.52 w=1 l=0.15
X11 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X12 Q a_713_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.1425 ps=1.285 w=1 l=0.15
X13 VGND D a_299_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X14 a_644_413# a_193_47# a_560_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0567 ps=0.69 w=0.42 l=0.15
X15 a_465_369# a_299_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.09575 pd=0.965 as=0.0864 ps=0.91 w=0.64 l=0.15
X16 a_560_47# a_27_47# a_465_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.09575 ps=0.965 w=0.42 l=0.15
X17 VGND GATE a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__decap_3 VPWR VGND VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
.ends

.subckt sky130_fd_sc_hd__buf_2 VPWR VGND VPB VNB X A
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o41a_4 VGND VPWR VPB VNB X B1 A4 A3 A2 A1
X0 a_467_47# A4 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_467_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.09425 pd=0.94 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VGND A1 a_467_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.15275 ps=1.12 w=0.65 l=0.15
X3 a_467_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.09425 pd=0.94 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_467_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.15275 pd=1.12 as=0.19825 ps=1.26 w=0.65 l=0.15
X5 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.135 ps=1.27 w=1 l=0.15
X6 VPWR A1 a_1083_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 a_1083_297# A2 a_889_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VGND A3 a_467_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 a_79_21# B1 a_467_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 a_889_297# A2 a_1083_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X13 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 a_639_297# A3 a_889_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X17 VGND A2 a_467_47# VNB sky130_fd_pr__nfet_01v8 ad=0.19825 pd=1.26 as=0.09425 ps=0.94 w=0.65 l=0.15
X18 a_889_297# A3 a_639_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 a_639_297# A4 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 VPWR B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.145 ps=1.29 w=1 l=0.15
X22 VGND A4 a_467_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.09425 ps=0.94 w=0.65 l=0.15
X23 a_1083_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.49 pd=2.98 as=0.135 ps=1.27 w=1 l=0.15
X24 a_79_21# A4 a_639_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X25 a_467_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.3185 pd=2.28 as=0.08775 ps=0.92 w=0.65 l=0.15
X26 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X27 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__decap_6 VPWR VGND VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
.ends

.subckt sky130_fd_sc_hd__or4_1 VPWR VGND VPB VNB B D C A X
X0 a_27_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_27_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_277_297# B a_205_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VPWR A a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.101875 ps=0.99 w=0.65 l=0.15
X5 a_205_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.14825 ps=1.34 w=1 l=0.15
X7 VGND C a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_109_297# D a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 VGND A a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__and2_1 VPWR VGND VPB VNB X A B
X0 VPWR B a_59_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 X a_59_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X2 VGND B a_145_75# VNB sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_59_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X4 X a_59_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X5 a_145_75# A a_59_75# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_2 VGND VPWR VPB VNB A X
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X1 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__dlymetal6s2s_1 VPWR VGND VPB VNB X A
X0 a_558_47# a_381_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X1 VGND X a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_841_47# a_664_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X3 VPWR A a_62_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 VGND A a_62_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 a_558_47# a_381_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X6 X a_62_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X7 VPWR X a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 a_841_47# a_664_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X9 X a_62_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X10 VPWR a_558_47# a_664_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X11 VGND a_558_47# a_664_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_4 VPWR VGND VPB VNB A X
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor2_1 VGND VPWR VPB VNB A B Y
X0 VPWR A a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_109_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VPWR VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
.ends

.subckt sky130_fd_sc_hd__dfrtp_1 VGND VPWR VPB VNB CLK D RESET_B Q
X0 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X3 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X4 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X5 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X7 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X10 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X12 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X13 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X14 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X15 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X16 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X18 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X19 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X20 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X21 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X22 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X23 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X24 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X25 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X26 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X27 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
.ends

.subckt sky130_fd_sc_hd__and2b_1 VGND VPWR VPB VNB A_N X B
X0 VPWR B a_207_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X1 X a_207_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X2 a_297_47# a_27_413# a_207_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 X a_207_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X4 a_207_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X5 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 VGND B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X7 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a22o_1 VPWR VGND VPB VNB B1 A1 A2 X B2
X0 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X1 a_27_297# B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X2 VGND A2 a_373_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X3 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X4 a_27_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X6 a_373_47# A1 a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X7 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X8 a_109_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 a_109_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and3_2 VPWR VGND VPB VNB X C B A
X0 VPWR a_29_311# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_29_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.15075 ps=1.345 w=1 l=0.15
X2 VPWR A a_29_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 VGND a_29_311# X VNB sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_184_53# B a_112_53# VNB sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X5 VPWR C a_29_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15075 pd=1.345 as=0.074375 ps=0.815 w=0.42 l=0.15
X6 X a_29_311# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1304 ps=1.105 w=0.65 l=0.15
X7 a_112_53# A a_29_311# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 a_29_311# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 VGND C a_184_53# VNB sky130_fd_pr__nfet_01v8 ad=0.1304 pd=1.105 as=0.05355 ps=0.675 w=0.42 l=0.15
.ends

.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
.ends

.subckt sky130_fd_sc_hd__nor4_2 VGND VPWR VPB VNB B D Y A C
X0 a_281_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_475_297# D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y D a_475_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VGND D Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X9 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 Y D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X12 a_475_297# C a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 a_281_297# C a_475_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X14 a_27_297# B a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X15 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__mux2_1 VGND VPWR VPB VNB X A1 S A0
X0 VPWR a_505_21# a_535_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1 a_505_21# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_218_374# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X3 VGND a_505_21# a_439_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_76_199# A0 a_218_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X5 a_505_21# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X6 a_439_47# A0 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X7 a_535_374# A1 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X8 a_76_199# A1 a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_218_47# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21o_1 VPWR VGND VPB VNB A2 A1 B1 X
X0 a_81_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X1 a_299_297# B1 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X2 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3 VPWR A1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X4 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X5 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X6 a_299_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7 a_384_47# A1 a_81_21# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4b_4 VGND VPWR VPB VNB X D_N C B A
X0 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 VGND a_215_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VPWR a_215_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_109_93# D_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10785 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 a_215_297# a_109_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.16535 ps=1.82 w=0.65 l=0.15
X5 VGND C a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1235 ps=1.03 w=0.65 l=0.15
X6 VGND A a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X8 a_215_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_109_93# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X10 VPWR A a_487_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.135 ps=1.27 w=1 l=0.15
X11 VGND a_215_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 a_487_297# B a_403_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 a_403_297# C a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X14 VPWR a_215_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X15 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1235 ps=1.03 w=0.65 l=0.15
X16 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 a_297_297# a_109_93# a_215_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a2111o_1 VGND VPWR VPB VNB A2 A1 B1 C1 D1 X
X0 VGND A2 a_660_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.082875 ps=0.905 w=0.65 l=0.15
X1 VGND C1 a_85_193# VNB sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.10075 ps=0.96 w=0.65 l=0.15
X2 a_414_297# C1 a_334_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X3 VGND a_85_193# X VNB sky130_fd_pr__nfet_01v8 ad=0.274625 pd=1.495 as=0.2145 ps=1.96 w=0.65 l=0.15
X4 a_334_297# D1 a_85_193# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X5 a_516_297# B1 a_414_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X6 a_516_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X7 a_660_47# A1 a_85_193# VNB sky130_fd_pr__nfet_01v8 ad=0.082875 pd=0.905 as=0.18525 ps=1.22 w=0.65 l=0.15
X8 a_85_193# D1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.274625 ps=1.495 w=0.65 l=0.15
X9 VPWR A1 a_516_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X10 a_85_193# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X11 VPWR a_85_193# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21a_1 VGND VPWR VPB VNB A1 A2 B1 X
X0 VPWR A1 a_382_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1525 ps=1.305 w=1 l=0.15
X1 a_297_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X2 a_297_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VGND A2 a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3275 pd=1.655 as=0.28 ps=2.56 w=1 l=0.15
X5 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.3275 ps=1.655 w=1 l=0.15
X6 a_382_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.195 ps=1.39 w=1 l=0.15
X7 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o221a_1 VGND VPWR VPB VNB B1 B2 A2 A1 X C1
X0 a_240_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1 X a_51_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VGND A1 a_240_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 a_51_297# B2 a_245_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.4125 pd=1.825 as=0.105 ps=1.21 w=1 l=0.15
X4 a_149_47# C1 a_51_297# VNB sky130_fd_pr__nfet_01v8 ad=0.099125 pd=0.955 as=0.2015 ps=1.92 w=0.65 l=0.15
X5 a_240_47# B1 a_149_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.099125 ps=0.955 w=0.65 l=0.15
X6 VPWR A1 a_512_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X7 X a_51_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.165 ps=1.33 w=1 l=0.15
X8 a_149_47# B2 a_240_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_245_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X10 VPWR C1 a_51_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.34 ps=2.68 w=1 l=0.15
X11 a_512_297# A2 a_51_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.4125 ps=1.825 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o22a_2 VGND VPWR VPB VNB A1 A2 B2 B1 X
X0 a_301_47# B2 a_81_21# VNB sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 VGND A2 a_301_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1235 ps=1.03 w=0.65 l=0.15
X2 a_383_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.39 ps=1.78 w=1 l=0.15
X3 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.39 pd=1.78 as=0.135 ps=1.27 w=1 l=0.15
X4 a_301_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 X a_81_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7 X a_81_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X8 VPWR A1 a_579_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.105 ps=1.21 w=1 l=0.15
X9 a_81_21# B1 a_301_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10 a_579_297# A2 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.235 ps=1.47 w=1 l=0.15
X11 a_81_21# B2 a_383_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.235 pd=1.47 as=0.105 ps=1.21 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__dlygate4sd3_1 VGND VPWR VPB VNB X A
X0 VPWR A a_49_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 VGND a_285_47# a_391_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.5
X2 X a_391_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X3 VGND A a_49_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 VPWR a_285_47# a_391_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.5
X5 a_285_47# a_49_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X6 a_285_47# a_49_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X7 X a_391_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a32o_1 VGND VPWR VPB VNB X A3 A2 A1 B1 B2
X0 a_93_21# A1 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.14625 ps=1.1 w=0.65 l=0.15
X1 a_93_21# B1 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X2 a_584_47# B1 a_93_21# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X3 VPWR a_93_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2425 pd=1.485 as=0.33 ps=2.66 w=1 l=0.15
X4 VGND B2 a_584_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.06825 ps=0.86 w=0.65 l=0.15
X5 a_256_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167375 ps=1.165 w=0.65 l=0.15
X6 a_250_297# B2 a_93_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7 VGND a_93_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.167375 pd=1.165 as=0.2145 ps=1.96 w=0.65 l=0.15
X8 a_250_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.2425 ps=1.485 w=1 l=0.15
X9 VPWR A2 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X10 a_250_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X11 a_346_47# A2 a_256_47# VNB sky130_fd_pr__nfet_01v8 ad=0.14625 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__diode_2 VGND VPWR VPB VNB DIODE
X0 VNB DIODE sky130_fd_pr__diode_pw2nd_05v5 perim=2.64e+06 area=4.347e+11
.ends

.subckt sky130_fd_sc_hd__dlygate4sd1_1 VPWR VGND VPB VNB X A
X0 X a_299_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X1 VPWR a_193_47# a_299_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5 VGND a_193_47# a_299_93# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 X a_299_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X7 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_4 VGND VPWR VPB VNB A X
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X6 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X8 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X9 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o211a_1 VGND VPWR VPB VNB X A1 A2 B1 C1
X0 VGND A1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1 a_510_47# B1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.143 ps=1.09 w=0.65 l=0.15
X2 a_79_21# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.175 ps=1.35 w=1 l=0.15
X3 VPWR B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.22 ps=1.44 w=1 l=0.15
X4 a_79_21# A2 a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.1625 ps=1.325 w=1 l=0.15
X5 a_297_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X6 a_79_21# C1 a_510_47# VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.11375 ps=1 w=0.65 l=0.15
X7 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X8 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X9 a_215_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.105625 ps=0.975 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__conb_1 VGND VPWR VPB VNB LO HI
X0 VPWR HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1 LO VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
.ends

.subckt sky130_fd_sc_hd__and4_1 VGND VPWR VPB VNB X D C B A
X0 a_27_47# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X1 a_197_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.31245 ps=1.68 w=1 l=0.15
X3 a_303_47# C a_197_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X4 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 VPWR D a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.31245 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X6 VGND D a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.196275 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X8 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196275 ps=1.33 w=0.65 l=0.15
X9 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand3b_1 VGND VPWR VPB VNB Y B C A_N
X0 Y a_53_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.1925 ps=1.385 w=1 l=0.15
X1 a_232_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X2 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1925 pd=1.385 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR A_N a_53_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 VGND A_N a_53_93# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 a_316_47# B a_232_47# VNB sky130_fd_pr__nfet_01v8 ad=0.125125 pd=1.035 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 Y a_53_93# a_316_47# VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.125125 ps=1.035 w=0.65 l=0.15
X7 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__dlymetal6s4s_1 VPWR VGND VPB VNB X A
X0 X a_345_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X1 VPWR a_239_47# a_345_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_841_47# a_664_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X3 VGND a_239_47# a_345_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 VPWR A a_62_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 VGND A a_62_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 X a_345_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X7 a_239_47# a_62_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X8 a_841_47# a_664_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X9 a_239_47# a_62_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X10 VPWR X a_664_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X11 VGND X a_664_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand2_1 VGND VPWR VPB VNB A Y B
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A a_113_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_113_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__decap_8 VPWR VGND VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
.ends

.subckt sky130_fd_sc_hd__and3_4 VGND VPWR VPB VNB X A B C
X0 VPWR A a_94_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1975 pd=1.395 as=0.305 ps=2.61 w=1 l=0.15
X1 a_294_47# B a_185_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.128375 ps=1.045 w=0.65 l=0.15
X2 a_185_47# A a_94_47# VNB sky130_fd_pr__nfet_01v8 ad=0.128375 pd=1.045 as=0.19825 ps=1.91 w=0.65 l=0.15
X3 VPWR a_94_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X4 VGND C a_294_47# VNB sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X5 a_94_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1975 ps=1.395 w=1 l=0.15
X6 X a_94_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X7 X a_94_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X8 VPWR C a_94_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X9 X a_94_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X10 VGND a_94_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X11 VPWR a_94_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 VGND a_94_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X13 X a_94_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a221o_1 VPWR VGND VPB VNB A1 A2 X B1 B2 C1
X0 a_465_47# A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X2 a_109_297# B1 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X5 a_205_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X6 VPWR A2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X7 a_193_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X8 a_27_47# B1 a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X9 a_109_297# C1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10 VGND C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X11 VGND A2 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3_1 VPWR VGND VPB VNB B C A X
X0 X a_29_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.14825 ps=1.34 w=1 l=0.15
X1 a_111_297# C a_29_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 X a_29_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.101875 ps=0.99 w=0.65 l=0.15
X3 a_183_297# B a_111_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 VPWR A a_183_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_29_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 VGND C a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7 VGND A a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand4_4 VPWR VGND VPB VNB C Y A B D
X0 a_27_47# C a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_27_47# C a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_445_47# B a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 a_445_47# B a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_27_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 a_27_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 Y A a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X14 Y A a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 a_803_47# B a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X17 a_803_47# B a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 VGND D a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 a_445_47# C a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 a_803_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X23 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X24 a_445_47# C a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X25 a_803_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X26 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X30 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X31 VGND D a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand2b_1 VGND VPWR VPB VNB A_N B Y
X0 VGND A_N a_27_93# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 Y a_27_93# a_206_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_206_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X3 VPWR a_27_93# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X4 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X5 VPWR A_N a_27_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__inv_2 VPWR VGND VPB VNB Y A
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21oi_1 VPWR VGND VPB VNB A2 A1 B1 Y
X0 a_199_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.095875 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X1 a_113_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1475 ps=1.295 w=1 l=0.15
X2 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X3 VPWR A1 a_113_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.14 ps=1.28 w=1 l=0.15
X4 a_113_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X5 VGND A2 a_199_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.095875 ps=0.945 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21ai_1 VGND VPWR VPB VNB A2 B1 Y A1
X0 Y A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X1 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X2 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X3 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X5 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o31a_1 VGND VPWR VPB VNB X A1 A2 A3 B1
X0 a_103_199# B1 a_253_47# VNB sky130_fd_pr__nfet_01v8 ad=0.2015 pd=1.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X1 VPWR a_103_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.36 ps=2.72 w=1 l=0.15
X2 a_337_297# A2 a_253_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3 a_103_199# A3 a_337_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2125 pd=1.425 as=0.165 ps=1.33 w=1 l=0.15
X4 a_253_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.195 ps=1.39 w=1 l=0.15
X5 VPWR B1 a_103_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.345 pd=2.69 as=0.2125 ps=1.425 w=1 l=0.15
X6 VGND a_103_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.234 ps=2.02 w=0.65 l=0.15
X7 a_253_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12675 ps=1.04 w=0.65 l=0.15
X8 a_253_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X9 VGND A2 a_253_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_1 VGND VPWR VPB VNB X A
X0 VPWR a_75_212# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1 a_75_212# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 a_75_212# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3 VGND a_75_212# X VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand3_1 VGND VPWR VPB VNB A B Y C
X0 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X2 a_193_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 Y A a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X4 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5 a_109_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and2_4 VGND VPWR VPB VNB A X B
X0 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X1 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X3 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 VGND B a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 a_110_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X7 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X8 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X9 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X10 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X11 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and3b_1 VGND VPWR VPB VNB B A_N X C
X0 a_109_93# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10785 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 X a_209_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X2 a_109_93# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1087 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 a_296_53# a_109_93# a_209_311# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.107825 ps=1.36 w=0.42 l=0.15
X4 VPWR C a_209_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.074375 ps=0.815 w=0.42 l=0.15
X5 a_368_53# B a_296_53# VNB sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 X a_209_311# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122275 ps=1.08 w=0.65 l=0.15
X7 a_209_311# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VPWR a_109_93# a_209_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1085 ps=1.36 w=0.42 l=0.15
X9 VGND C a_368_53# VNB sky130_fd_pr__nfet_01v8 ad=0.122275 pd=1.08 as=0.05355 ps=0.675 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand2_4 VGND VPWR VPB VNB B Y A
X0 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a211o_1 VGND VPWR VPB VNB X C1 A2 A1 B1
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X1 a_80_21# C1 a_472_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X2 VPWR A2 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.17225 ps=1.83 w=0.65 l=0.15
X5 a_300_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X6 a_217_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7 a_80_21# A1 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X8 a_472_297# B1 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X9 a_80_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o22a_1 VGND VPWR VPB VNB B2 A2 A1 B1 X
X0 a_78_199# B1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1 VPWR A1 a_493_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2 a_493_297# A2 a_78_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.235 ps=1.47 w=1 l=0.15
X3 VPWR a_78_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3725 pd=1.745 as=0.28 ps=2.56 w=1 l=0.15
X4 VGND A2 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.11375 ps=1 w=0.65 l=0.15
X5 a_78_199# B2 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.235 pd=1.47 as=0.1175 ps=1.235 w=1 l=0.15
X6 a_215_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 a_215_47# B2 a_78_199# VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 a_292_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1175 pd=1.235 as=0.3725 ps=1.745 w=1 l=0.15
X9 VGND a_78_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand2b_2 VGND VPWR VPB VNB A_N Y B
X0 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.335 ps=1.67 w=1 l=0.15
X1 VGND A_N a_27_93# VNB sky130_fd_pr__nfet_01v8 ad=0.194 pd=1.95 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 VGND B a_229_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 Y a_27_93# a_229_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4 a_229_47# a_27_93# Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y a_27_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.1468 ps=1.34 w=1 l=0.15
X6 VPWR a_27_93# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.335 pd=1.67 as=0.165 ps=1.33 w=1 l=0.15
X7 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.135 ps=1.27 w=1 l=0.15
X8 a_229_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VPWR A_N a_27_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1468 pd=1.34 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__mux4_1 VGND VPWR VPB VNB A1 A0 S0 A3 A2 S1 X
X0 a_277_47# a_247_21# a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 VGND S0 a_247_21# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_834_97# a_247_21# a_750_97# VNB sky130_fd_pr__nfet_01v8 ad=0.10795 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 VGND A3 a_668_97# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1079 ps=1.36 w=0.42 l=0.15
X4 a_1290_413# S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 a_834_97# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 a_750_97# S0 a_757_363# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1079 ps=1.36 w=0.42 l=0.15
X7 a_27_47# S0 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.085225 ps=0.925 w=0.42 l=0.15
X8 X a_1478_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X9 VPWR A1 a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10 VPWR S0 a_247_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1079 pd=1.36 as=0.1083 ps=1.36 w=0.42 l=0.15
X11 X a_1478_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X12 a_193_47# A0 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 a_750_97# a_1290_413# a_1478_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2688 pd=2.12 as=0.092075 ps=0.99 w=0.42 l=0.15
X14 a_1478_413# S1 a_277_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.092075 pd=0.99 as=0.1092 ps=1.36 w=0.42 l=0.15
X15 a_1290_413# S1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X16 a_277_47# a_247_21# a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0.085225 pd=0.925 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 a_750_97# S0 a_668_97# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X18 a_923_363# a_247_21# a_750_97# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.090125 pd=0.995 as=0.0567 ps=0.69 w=0.42 l=0.15
X19 a_757_363# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X20 VPWR A3 a_923_363# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.090125 ps=0.995 w=0.42 l=0.15
X21 a_277_47# a_1290_413# a_1478_413# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.151025 ps=1.285 w=0.42 l=0.15
X22 a_193_413# A0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X23 a_193_413# S0 a_277_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1079 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X24 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X25 a_1478_413# S1 a_750_97# VNB sky130_fd_pr__nfet_01v8 ad=0.151025 pd=1.285 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4_4 VPWR VGND VPB VNB D C B A X
X0 VPWR A a_304_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.135 ps=1.27 w=1 l=0.15
X1 a_304_297# B a_220_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND C a_32_297# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1235 ps=1.03 w=0.65 l=0.15
X3 a_220_297# C a_114_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X4 a_32_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.169 ps=1.82 w=0.65 l=0.15
X5 a_32_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VPWR a_32_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X7 X a_32_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VGND A a_32_297# VNB sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VPWR a_32_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 X a_32_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1235 ps=1.03 w=0.65 l=0.15
X11 X a_32_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 X a_32_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X13 a_114_297# D a_32_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.26 ps=2.52 w=1 l=0.15
X14 VGND a_32_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 VGND a_32_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a31o_1 VGND VPWR VPB VNB X A3 A2 A1 B1
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X1 a_209_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X2 a_303_47# A2 a_209_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X3 a_209_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X5 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X6 a_80_21# A1 a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X7 VPWR A2 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X8 a_80_21# B1 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X9 a_209_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__or2_1 VGND VPWR VPB VNB X A B
X0 VGND A a_68_297# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_68_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 X a_68_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X3 VPWR A a_150_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 X a_68_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X5 a_150_297# B a_68_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o211a_4 VGND VPWR VPB VNB X C1 B1 A2 A1
X0 VGND A1 a_474_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.104 ps=0.97 w=0.65 l=0.15
X1 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 VPWR A1 a_1122_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2525 pd=1.505 as=0.14 ps=1.28 w=1 l=0.15
X5 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.19175 pd=1.89 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VPWR C1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.2525 ps=1.505 w=1 l=0.15
X8 a_950_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.16 ps=1.32 w=1 l=0.15
X9 a_557_47# B1 a_474_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X10 a_474_47# B1 a_748_47# VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.091 ps=0.93 w=0.65 l=0.15
X11 VGND A2 a_474_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X12 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 a_79_21# C1 a_557_47# VNB sky130_fd_pr__nfet_01v8 ad=0.144625 pd=1.095 as=0.06825 ps=0.86 w=0.65 l=0.15
X15 a_474_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X16 a_79_21# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.14 ps=1.28 w=1 l=0.15
X17 a_748_47# C1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.144625 ps=1.095 w=0.65 l=0.15
X18 a_474_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.12675 ps=1.04 w=0.65 l=0.15
X19 VPWR B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.195 ps=1.39 w=1 l=0.15
X20 a_79_21# A2 a_950_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X21 a_1122_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X22 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X23 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__xnor2_1 VGND VPWR VPB VNB B A Y
X0 a_377_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.365 ps=1.73 w=1 l=0.15
X1 a_47_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3 ps=2.6 w=1 l=0.15
X2 a_129_47# B a_47_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_285_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4 Y a_47_47# a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VGND A a_129_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.06825 ps=0.86 w=0.65 l=0.15
X6 VPWR A a_47_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.365 pd=1.73 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR a_47_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.165 ps=1.33 w=1 l=0.15
X8 Y B a_377_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o211a_2 VPWR VGND VPB VNB A2 A1 X C1 B1
X0 a_27_47# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3675 pd=1.735 as=0.14 ps=1.28 w=1 l=0.15
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.23075 pd=2.01 as=0.091 ps=0.93 w=0.65 l=0.15
X2 VPWR C1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3 VPWR A1 a_373_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X4 a_182_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.16535 ps=1.82 w=0.65 l=0.15
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.195 ps=1.39 w=1 l=0.15
X6 a_182_47# B1 a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.16535 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.104 ps=0.97 w=0.65 l=0.15
X8 a_373_297# A2 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.3675 ps=1.735 w=1 l=0.15
X9 a_110_47# C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X10 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X11 VGND A1 a_182_47# VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3b_1 VGND VPWR VPB VNB B C_N A X
X0 a_109_93# C_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 a_215_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 VGND a_109_93# a_215_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 VGND A a_215_53# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 VPWR A a_369_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06825 ps=0.745 w=0.42 l=0.15
X5 a_369_297# B a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 X a_215_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X7 a_297_297# a_109_93# a_215_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 a_109_93# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 X a_215_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.10025 ps=0.985 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a22oi_1 VPWR VGND VPB VNB B2 B1 Y A1 A2
X0 Y B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X1 Y B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.135 ps=1.27 w=1 l=0.15
X3 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 a_381_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X5 a_109_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 a_109_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X7 VGND A2 a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.234 pd=2.02 as=0.06825 ps=0.86 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_8 VGND VPWR VPB VNB X A
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.1134 pd=1.38 as=0.0588 ps=0.7 w=0.42 l=0.15
X10 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X11 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X14 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X16 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X17 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X18 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X19 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a2111oi_2 VGND VPWR VPB VNB A1 A2 D1 C1 B1 Y
X0 a_467_297# B1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.16 ps=1.32 w=1 l=0.15
X1 a_287_297# D1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 VPWR A2 a_467_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.14 ps=1.28 w=1 l=0.15
X3 a_923_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.112125 ps=0.995 w=0.65 l=0.15
X4 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.12675 ps=1.04 w=0.65 l=0.15
X5 a_28_297# B1 a_467_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14 ps=1.28 w=1 l=0.15
X6 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.18525 ps=1.87 w=0.65 l=0.15
X7 a_28_297# C1 a_287_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.14 ps=1.28 w=1 l=0.15
X8 Y A1 a_923_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X9 VGND A2 a_684_47# VNB sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17875 ps=1.2 w=0.65 l=0.15
X10 Y D1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X11 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.105625 ps=0.975 w=0.65 l=0.15
X12 Y D1 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13 a_467_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.335 pd=2.67 as=0.16 ps=1.32 w=1 l=0.15
X14 VGND D1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.091 ps=0.93 w=0.65 l=0.15
X15 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.12675 ps=1.04 w=0.65 l=0.15
X16 VPWR A1 a_467_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.26 ps=2.52 w=1 l=0.15
X17 a_115_297# C1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.285 ps=2.57 w=1 l=0.15
X18 a_467_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X19 a_684_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.2 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__inv_8 VGND VPWR VPB VNB Y A
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfrtp_4 VGND VPWR VPB VNB CLK D RESET_B Q
X0 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X3 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X4 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X5 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X12 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X14 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X15 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X16 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X17 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X18 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X19 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X20 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X21 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X22 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X23 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X24 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X25 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X26 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X27 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X28 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X29 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X30 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X31 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X32 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X33 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21ba_1 VGND VPWR VPB VNB B1_N A1 A2 X
X0 a_222_93# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X1 VPWR A1 a_544_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.105 ps=1.21 w=1 l=0.15
X2 VGND a_79_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_222_93# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.18575 ps=1.415 w=0.42 l=0.15
X4 VGND A2 a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X5 a_448_47# a_222_93# a_79_199# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X6 a_79_199# a_222_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.3 ps=2.6 w=1 l=0.15
X7 a_544_297# A2 a_79_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X8 a_448_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VPWR a_79_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18575 pd=1.415 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o22a_4 VGND VPWR VPB VNB A1 B1 B2 A2 X
X0 VPWR B1 a_566_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X1 a_484_47# B1 a_96_21# VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 X a_96_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VPWR a_96_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_96_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 a_566_297# B2 a_96_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VPWR a_96_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 X a_96_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X8 VGND a_96_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_96_21# B2 a_566_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR A1 a_918_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.135 ps=1.27 w=1 l=0.15
X11 a_484_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 a_566_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X13 a_484_47# B2 a_96_21# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 a_96_21# A2 a_918_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 a_918_297# A2 a_96_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 a_484_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 a_918_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X18 a_96_21# B1 a_484_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X19 VGND A2 a_484_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 a_96_21# B2 a_484_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 VGND A1 a_484_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.11375 ps=1 w=0.65 l=0.15
X22 X a_96_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X23 VGND a_96_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__dlxtn_1 VGND VPWR VPB VNB Q D GATE_N
X0 VPWR D a_299_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1 a_560_47# a_27_47# a_465_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.054 pd=0.66 as=0.066 ps=0.745 w=0.36 l=0.15
X2 a_465_47# a_299_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 VPWR GATE_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4 VGND a_560_47# a_715_21# VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X5 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 VPWR a_560_47# a_715_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X7 a_650_47# a_193_47# a_560_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.054 ps=0.66 w=0.36 l=0.15
X8 Q a_715_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X9 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10 VPWR a_715_21# a_644_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07455 ps=0.775 w=0.42 l=0.15
X11 VGND D a_299_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X12 Q a_715_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X13 a_644_413# a_27_47# a_560_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07455 pd=0.775 as=0.0567 ps=0.69 w=0.42 l=0.15
X14 a_465_369# a_299_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.09575 pd=0.965 as=0.0864 ps=0.91 w=0.64 l=0.15
X15 a_560_47# a_193_47# a_465_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.09575 ps=0.965 w=0.42 l=0.15
X16 VGND GATE_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X17 VGND a_715_21# a_650_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor3b_2 VGND VPWR VPB VNB A Y C_N B
X0 a_281_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND a_531_21# Y VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 VPWR C_N a_531_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X7 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X9 a_281_297# a_531_21# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X10 Y a_531_21# a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X11 VGND C_N a_531_21# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X12 a_27_297# B a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X13 Y a_531_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__inv_16 VGND VPWR VPB VNB Y A
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X17 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X22 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X26 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X28 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X29 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X30 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X31 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o32a_4 VGND VPWR VPB VNB A2 A3 B2 X A1 B1
X0 a_27_47# B2 a_549_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 VGND a_549_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VPWR a_549_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 a_27_297# A2 a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4 a_277_297# A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 a_549_297# B2 a_739_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.135 ps=1.27 w=1 l=0.15
X6 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 a_739_297# B2 a_549_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15 ps=1.3 w=1 l=0.15
X9 a_739_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.09425 pd=0.94 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 a_549_297# B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0975 ps=0.95 w=0.65 l=0.15
X13 a_277_297# A3 a_549_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X14 VPWR B1 a_739_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15 X a_549_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 a_27_47# B1 a_549_297# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X17 a_549_297# A3 a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X18 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.09425 ps=0.94 w=0.65 l=0.15
X19 VPWR a_549_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VGND a_549_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 X a_549_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X23 a_549_297# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X24 X a_549_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X25 X a_549_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X26 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X27 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or2_2 VPWR VGND VPB VNB X A B
X0 a_121_297# B a_39_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 X a_39_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10675 ps=1.005 w=0.65 l=0.15
X2 VPWR a_39_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 X a_39_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.15575 ps=1.355 w=1 l=0.15
X4 VGND a_39_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VPWR A a_121_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15575 pd=1.355 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 VGND A a_39_297# VNB sky130_fd_pr__nfet_01v8 ad=0.10675 pd=1.005 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 a_39_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o311a_1 VGND VPWR VPB VNB X A1 A2 A3 B1 C1
X0 a_585_47# B1 a_266_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.118625 ps=1.015 w=0.65 l=0.15
X1 VGND A2 a_266_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1365 pd=1.07 as=0.117 ps=1.01 w=0.65 l=0.15
X2 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3125 pd=1.625 as=0.26 ps=2.52 w=1 l=0.15
X3 a_81_21# C1 a_585_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X4 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.203125 pd=1.275 as=0.169 ps=1.82 w=0.65 l=0.15
X5 a_266_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.3125 ps=1.625 w=1 l=0.15
X6 a_368_297# A2 a_266_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.18 ps=1.36 w=1 l=0.15
X7 a_266_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.118625 pd=1.015 as=0.1365 ps=1.07 w=0.65 l=0.15
X8 a_266_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.203125 ps=1.275 w=0.65 l=0.15
X9 a_81_21# A3 a_368_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.21 ps=1.42 w=1 l=0.15
X10 a_81_21# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15 ps=1.3 w=1 l=0.15
X11 VPWR B1 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.1375 ps=1.275 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o32a_1 VPWR VGND VPB VNB X A1 A2 A3 B2 B1
X0 a_77_199# B2 a_227_47# VNB sky130_fd_pr__nfet_01v8 ad=0.13325 pd=1.06 as=0.12675 ps=1.04 w=0.65 l=0.15
X1 a_323_297# A2 a_227_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.165 ps=1.33 w=1 l=0.15
X2 a_227_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3 a_227_47# B1 a_77_199# VNB sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.13325 ps=1.06 w=0.65 l=0.15
X4 VGND a_77_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5 VPWR B1 a_539_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.205 ps=1.41 w=1 l=0.15
X6 a_227_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X7 VPWR a_77_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.335 ps=2.67 w=1 l=0.15
X8 a_77_199# A3 a_323_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X9 VGND A2 a_227_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.10725 ps=0.98 w=0.65 l=0.15
X10 a_227_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 a_539_297# B2 a_77_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=1.41 as=0.195 ps=1.39 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_6 VPWR VGND VPB VNB A X
X0 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_161_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND A a_161_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 VPWR A a_161_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 a_161_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor3b_1 VGND VPWR VPB VNB C_N B Y A
X0 VGND a_91_199# Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.221 ps=1.98 w=0.65 l=0.15
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VPWR A a_245_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X3 a_91_199# C_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 a_245_297# B a_161_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_91_199# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X7 a_161_297# a_91_199# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.32 ps=2.64 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__inv_12 VGND VPWR VPB VNB Y A
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.515 pd=3.03 as=0.135 ps=1.27 w=1 l=0.15
X4 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.33475 pd=2.33 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X14 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o2bb2a_1 VPWR VGND VPB VNB X A1_N A2_N B2 B1
X0 a_206_369# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.14575 ps=1.335 w=0.42 l=0.15
X1 a_206_369# A2_N a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06615 ps=0.735 w=0.42 l=0.15
X2 VGND B2 a_489_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_585_369# B2 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0672 ps=0.74 w=0.42 l=0.15
X4 a_489_47# a_206_369# a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 a_489_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 VPWR A2_N a_206_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.20925 pd=1.345 as=0.129 ps=1.18 w=0.42 l=0.15
X7 a_76_199# a_206_369# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.20925 ps=1.345 w=0.42 l=0.15
X8 a_205_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06615 pd=0.735 as=0.098625 ps=0.98 w=0.42 l=0.15
X9 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.26 ps=2.52 w=1 l=0.15
X10 VPWR B1 a_585_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.098625 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3b_4 VGND VPWR VPB VNB C_N X A B
X0 a_176_21# a_27_47# a_626_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X1 a_626_297# B a_542_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR C_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 VGND a_176_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_542_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR a_176_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 X a_176_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 X a_176_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X8 X a_176_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_176_21# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 VPWR a_176_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 X a_176_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X12 a_176_21# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X13 VGND a_176_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 VGND B a_176_21# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 VGND C_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_1 VGND VPWR VPB VNB X A
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkinv_8 VGND VPWR VPB VNB A Y
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.135 ps=1.27 w=1 l=0.15
X6 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1375 ps=1.275 w=1 l=0.15
X11 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X16 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X19 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o41a_2 VGND VPWR VPB VNB A1 A2 A3 A4 B1 X
X0 VGND A2 a_393_47# VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.11375 ps=1 w=0.65 l=0.15
X1 a_496_297# A4 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.3025 ps=1.605 w=1 l=0.15
X2 a_393_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.115375 ps=1.005 w=0.65 l=0.15
X3 VPWR A1 a_697_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.41 pd=2.82 as=0.175 ps=1.35 w=1 l=0.15
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3025 pd=1.605 as=0.305 ps=1.61 w=1 l=0.15
X7 VGND A4 a_393_47# VNB sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.118625 ps=1.015 w=0.65 l=0.15
X8 a_697_297# A2 a_597_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.175 ps=1.35 w=1 l=0.15
X9 a_393_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.2665 pd=2.12 as=0.11375 ps=1 w=0.65 l=0.15
X10 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11 a_393_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.118625 pd=1.015 as=0.208 ps=1.94 w=0.65 l=0.15
X12 a_597_297# A3 a_496_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.1775 ps=1.355 w=1 l=0.15
X13 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_16 VGND VPWR VPB VNB A X
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X6 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X7 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X14 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X16 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X17 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X18 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X19 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X20 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X21 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X22 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X23 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X24 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X25 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X26 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X27 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X28 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X29 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X30 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X31 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X32 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X33 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X34 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X35 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X36 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X37 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X38 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X39 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21bo_1 VGND VPWR VPB VNB X A2 A1 B1_N
X0 a_298_297# a_27_413# a_215_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1 a_215_297# a_27_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1359 ps=1.1 w=0.65 l=0.15
X2 a_298_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.258375 ps=1.445 w=0.65 l=0.15
X4 VPWR B1_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X6 a_382_47# A1 a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VGND B1_N a_27_413# VNB sky130_fd_pr__nfet_01v8 ad=0.1359 pd=1.1 as=0.1113 ps=1.37 w=0.42 l=0.15
X8 VPWR A1 a_298_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X9 VGND A2 a_382_47# VNB sky130_fd_pr__nfet_01v8 ad=0.258375 pd=1.445 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkinv_4 VPWR VGND VPB VNB A Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.1659 pd=1.63 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.345 pd=2.69 as=0.14 ps=1.28 w=1 l=0.15
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.305 ps=2.61 w=1 l=0.15
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1386 ps=1.5 w=0.42 l=0.15
X8 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a22oi_2 VPWR VGND VPB VNB B2 B1 Y A1 A2
X0 a_109_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_467_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_467_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 Y B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 Y A1 a_467_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6 a_109_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND A2 a_467_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 Y B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_27_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 VPWR A1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 a_109_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15 VGND B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__xor2_1 VPWR VGND VPB VNB A X B
X0 X a_35_297# a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X1 X B a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_35_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_117_297# B a_35_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 VPWR B a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND A a_35_297# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25025 ps=1.42 w=0.65 l=0.15
X7 a_285_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR A a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__bufinv_16 VGND VPWR VPB VNB A Y
X0 a_361_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 VPWR a_361_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_361_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 Y a_361_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 VPWR a_361_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 Y a_361_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 Y a_361_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR a_27_47# a_361_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR a_361_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9 VPWR a_361_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VGND a_361_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 a_361_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 VGND a_361_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 VGND a_361_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 VGND a_361_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 VGND a_361_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 Y a_361_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 VGND a_361_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 VPWR a_361_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 Y a_361_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X22 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X23 a_361_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X24 Y a_361_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 Y a_361_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X26 VPWR a_27_47# a_361_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 Y a_361_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X28 Y a_361_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 Y a_361_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X30 a_361_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X31 VPWR a_361_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X32 Y a_361_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X33 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X34 VGND a_27_47# a_361_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X35 VPWR a_27_47# a_361_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X36 Y a_361_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X37 VGND a_27_47# a_361_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X38 VGND a_27_47# a_361_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X39 a_361_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X40 VPWR a_361_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X41 VPWR a_361_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X42 VGND a_361_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X43 VGND a_361_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X44 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X45 Y a_361_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X46 Y a_361_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X47 Y a_361_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X48 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X49 Y a_361_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a311o_1 VGND VPWR VPB VNB C1 B1 A1 A2 A3 X
X0 a_75_199# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.134875 ps=1.065 w=0.65 l=0.15
X1 a_208_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.125125 pd=1.035 as=0.112125 ps=0.995 w=0.65 l=0.15
X2 a_315_47# A2 a_208_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.17 as=0.125125 ps=1.035 w=0.65 l=0.15
X3 VGND B1 a_75_199# VNB sky130_fd_pr__nfet_01v8 ad=0.134875 pd=1.065 as=0.105625 ps=0.975 w=0.65 l=0.15
X4 a_75_199# A1 a_315_47# VNB sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.169 ps=1.17 w=0.65 l=0.15
X5 a_75_199# C1 a_544_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2075 ps=1.415 w=1 l=0.15
X6 a_544_297# B1 a_201_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2075 pd=1.415 as=0.1625 ps=1.325 w=1 l=0.15
X7 VPWR a_75_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1425 pd=1.285 as=0.285 ps=2.57 w=1 l=0.15
X8 a_201_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.1425 ps=1.285 w=1 l=0.15
X9 VPWR A2 a_201_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.165 ps=1.33 w=1 l=0.15
X10 a_201_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.305 ps=1.61 w=1 l=0.15
X11 VGND a_75_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o22ai_1 VGND VPWR VPB VNB A1 A2 B1 B2 Y
X0 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X1 a_27_47# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.092625 ps=0.935 w=0.65 l=0.15
X2 VPWR A1 a_307_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.105 ps=1.21 w=1 l=0.15
X3 a_307_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.2325 ps=1.465 w=1 l=0.15
X4 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2325 pd=1.465 as=0.1125 ps=1.225 w=1 l=0.15
X6 a_109_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1125 pd=1.225 as=0.26 ps=2.52 w=1 l=0.15
X7 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.092625 pd=0.935 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a2111oi_1 VPWR VGND VPB VNB D1 C1 B1 A1 Y A2
X0 a_316_297# C1 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.1725 ps=1.345 w=1 l=0.15
X1 Y D1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.125125 pd=1.035 as=0.481 ps=2.78 w=0.65 l=0.15
X2 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.12025 pd=1.02 as=0.125125 ps=1.035 w=0.65 l=0.15
X3 a_420_297# B1 a_316_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=1.58 as=0.185 ps=1.37 w=1 l=0.15
X4 VPWR A1 a_420_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.29 ps=1.58 w=1 l=0.15
X5 VGND A2 a_568_47# VNB sky130_fd_pr__nfet_01v8 ad=0.19175 pd=1.89 as=0.0845 ps=0.91 w=0.65 l=0.15
X6 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.19175 pd=1.24 as=0.12025 ps=1.02 w=0.65 l=0.15
X7 a_420_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.1375 ps=1.275 w=1 l=0.15
X8 a_217_297# D1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.755 ps=3.51 w=1 l=0.15
X9 a_568_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0845 pd=0.91 as=0.19175 ps=1.24 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__inv_6 VPWR VGND VPB VNB Y A
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.247 ps=2.06 w=0.65 l=0.15
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.43 ps=2.86 w=1 l=0.15
X9 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a2bb2o_1 VGND VPWR VPB VNB B1 B2 A2_N A1_N X
X0 a_226_47# A2_N a_226_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0441 ps=0.63 w=0.42 l=0.15
X1 a_489_413# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 a_226_297# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.16675 ps=1.435 w=0.42 l=0.15
X3 VPWR B2 a_489_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 a_489_413# a_226_47# a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 a_76_199# a_226_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1386 ps=1.08 w=0.42 l=0.15
X6 VGND B1 a_556_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 a_556_47# B2 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VGND A2_N a_226_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1386 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 a_226_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1201 ps=1.085 w=0.42 l=0.15
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16675 pd=1.435 as=0.26 ps=2.52 w=1 l=0.15
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.1201 pd=1.085 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfxtp_1 VPWR VGND VPB VNB CLK D Q
X0 Q a_1059_315# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_891_413# a_193_47# a_634_159# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2 a_561_413# a_27_47# a_466_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X3 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4 Q a_1059_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 VGND a_634_159# a_592_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X7 VPWR a_891_413# a_1059_315# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X8 a_466_413# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X9 VPWR a_634_159# a_561_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X10 a_634_159# a_466_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X11 a_634_159# a_466_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X12 a_975_413# a_193_47# a_891_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 VGND a_1059_315# a_1017_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X14 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X15 a_891_413# a_27_47# a_634_159# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X16 a_592_47# a_193_47# a_466_413# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X17 VPWR a_1059_315# a_975_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X18 a_1017_47# a_27_47# a_891_413# VNB sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X19 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X20 a_466_413# a_27_47# a_381_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X21 VGND a_891_413# a_1059_315# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X22 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X23 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__and4b_1 VGND VPWR VPB VNB X D C B A_N
X0 a_297_47# a_27_47# a_193_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 a_369_47# B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0441 ps=0.63 w=0.42 l=0.15
X2 VPWR D a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.06615 ps=0.735 w=0.42 l=0.15
X3 X a_193_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1034 ps=1 w=0.65 l=0.15
X4 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 VGND D a_469_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1034 pd=1 as=0.0609 ps=0.71 w=0.42 l=0.15
X6 X a_193_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X7 VPWR B a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1281 pd=1.03 as=0.0987 ps=0.89 w=0.42 l=0.15
X8 a_193_413# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.1281 ps=1.03 w=0.42 l=0.15
X9 a_193_413# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 a_469_47# C a_369_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0735 ps=0.77 w=0.42 l=0.15
X11 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkinv_16 VGND VPWR VPB VNB Y A
X0 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.14 ps=1.28 w=1 l=0.15
X3 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.2175 ps=1.435 w=1 l=0.15
X13 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.06615 pd=0.735 as=0.0588 ps=0.7 w=0.42 l=0.15
X14 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.275 ps=2.55 w=1 l=0.15
X15 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X16 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X17 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X18 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X19 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X20 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X21 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X22 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X23 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X24 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2175 pd=1.435 as=0.1575 ps=1.315 w=1 l=0.15
X25 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X26 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X27 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X28 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X29 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X30 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X31 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X32 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X33 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X34 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.09135 pd=0.855 as=0.06615 ps=0.735 w=0.42 l=0.15
X35 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X36 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X37 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X38 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X39 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.09135 ps=0.855 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor4_1 VGND VPWR VPB VNB Y D C B A
X0 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.089375 ps=0.925 w=0.65 l=0.15
X1 a_191_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.13 ps=1.26 w=1 l=0.15
X2 VPWR A a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.118625 ps=1.015 w=0.65 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 a_297_297# B a_191_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X6 a_109_297# D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.13 pd=1.26 as=0.26 ps=2.52 w=1 l=0.15
X7 Y D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.118625 pd=1.015 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4b_1 VPWR VGND VPB VNB B C A X D_N
X0 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X1 a_109_53# D_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_215_297# a_109_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.101875 ps=0.99 w=0.65 l=0.15
X4 a_392_297# C a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.04515 pd=0.635 as=0.06825 ps=0.745 w=0.42 l=0.15
X5 a_465_297# B a_392_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06405 pd=0.725 as=0.04515 ps=0.635 w=0.42 l=0.15
X6 a_215_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 VPWR A a_465_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06405 ps=0.725 w=0.42 l=0.15
X8 a_297_297# a_109_53# a_215_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 a_109_53# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X10 VGND C a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06405 ps=0.725 w=0.42 l=0.15
X11 VGND A a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__or2_4 VGND VPWR VPB VNB B A X
X0 a_121_297# B a_35_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X1 VPWR a_35_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X2 X a_35_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 X a_35_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X4 X a_35_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VPWR a_35_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 X a_35_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X7 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VPWR A a_121_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X9 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 VGND A a_35_297# VNB sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 a_35_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o2111a_1 VPWR VGND VPB VNB X D1 C1 B1 A2 A1
X0 a_676_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.2125 ps=1.425 w=1 l=0.15
X1 a_512_47# B1 a_409_47# VNB sky130_fd_pr__nfet_01v8 ad=0.19825 pd=1.26 as=0.118625 ps=1.015 w=0.65 l=0.15
X2 a_306_47# D1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.118625 pd=1.015 as=0.19825 ps=1.91 w=0.65 l=0.15
X3 VGND A2 a_512_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.19825 ps=1.26 w=0.65 l=0.15
X4 VPWR C1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.2175 ps=1.435 w=1 l=0.15
X5 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2125 pd=1.425 as=0.305 ps=1.61 w=1 l=0.15
X6 VPWR A1 a_676_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.105 ps=1.21 w=1 l=0.15
X7 a_512_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 a_409_47# C1 a_306_47# VNB sky130_fd_pr__nfet_01v8 ad=0.118625 pd=1.015 as=0.118625 ps=1.015 w=0.65 l=0.15
X9 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3825 pd=1.765 as=0.26 ps=2.52 w=1 l=0.15
X10 a_79_21# D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2175 pd=1.435 as=0.3825 ps=1.765 w=1 l=0.15
X11 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o32ai_4 VGND VPWR VPB VNB B2 Y B1 A3 A2 A1
X0 a_1224_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 VPWR A1 a_1224_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1825 ps=1.365 w=1 l=0.15
X2 a_27_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1425 pd=1.285 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_806_297# A3 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.20475 ps=1.28 w=0.65 l=0.15
X8 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.20475 pd=1.28 as=0.13975 ps=1.08 w=0.65 l=0.15
X10 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_806_297# A3 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 Y A3 a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 a_27_47# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 a_27_47# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0.092625 pd=0.935 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 Y A3 a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X19 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.118625 ps=1.015 w=0.65 l=0.15
X22 a_27_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.092625 ps=0.935 w=0.65 l=0.15
X24 a_806_297# A2 a_1224_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X25 Y B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X26 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X27 VPWR B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1425 ps=1.285 w=1 l=0.15
X28 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X29 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.13975 pd=1.08 as=0.08775 ps=0.92 w=0.65 l=0.15
X30 a_1224_297# A2 a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X31 a_1224_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.135 ps=1.27 w=1 l=0.15
X32 a_806_297# A2 a_1224_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X33 VPWR A1 a_1224_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X34 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X35 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X36 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25675 ps=1.44 w=0.65 l=0.15
X37 a_1224_297# A2 a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X38 Y B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X39 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.118625 pd=1.015 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor2_2 VGND VPWR VPB VNB B Y A
X0 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X5 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X7 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o211ai_1 VGND VPWR VPB VNB A1 Y C1 B1 A2
X0 a_110_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.265 ps=2.53 w=1 l=0.15
X1 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.17225 ps=1.83 w=0.65 l=0.15
X2 Y A2 a_110_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X3 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X4 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X5 a_326_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.12675 ps=1.04 w=0.65 l=0.15
X6 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.635 pd=3.27 as=0.195 ps=1.39 w=1 l=0.15
X7 Y C1 a_326_47# VNB sky130_fd_pr__nfet_01v8 ad=0.39325 pd=2.51 as=0.06825 ps=0.86 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o41ai_2 VGND VPWR VPB VNB A1 A2 A3 A4 Y B1
X0 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 VGND A4 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X4 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 a_299_297# A3 a_549_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X9 a_549_297# A3 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 a_299_297# A4 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 Y A4 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12 a_743_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X13 VPWR A1 a_743_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 a_743_297# A2 a_549_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 a_27_47# A4 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X16 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X17 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 a_549_297# A2 a_743_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X19 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a221o_2 VPWR VGND VPB VNB C1 B2 B1 A1 A2 X
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.135 ps=1.27 w=1 l=0.15
X1 a_465_47# A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1575 ps=1.315 w=1 l=0.15
X3 a_109_297# B1 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.102375 ps=0.965 w=0.65 l=0.15
X6 a_205_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X7 VPWR A2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X8 a_193_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X9 a_27_47# B1 a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X10 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 a_109_297# C1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12 VGND C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X13 VGND A2 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a31oi_1 VGND VPWR VPB VNB A3 A2 A1 Y B1
X0 Y A1 a_181_47# VNB sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.118625 ps=1.015 w=0.65 l=0.15
X1 a_181_47# A2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.118625 pd=1.015 as=0.06825 ps=0.86 w=0.65 l=0.15
X2 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.105625 ps=0.975 w=0.65 l=0.15
X3 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.135 ps=1.27 w=1 l=0.15
X4 Y B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1625 ps=1.325 w=1 l=0.15
X5 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.1525 ps=1.305 w=1 l=0.15
X6 a_109_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 a_109_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o221ai_4 VGND VPWR VPB VNB B2 Y A2 A1 B1 C1
X0 a_471_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_471_47# B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_471_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR A1 a_1241_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.295 pd=2.59 as=0.135 ps=1.27 w=1 l=0.15
X5 a_471_47# B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_471_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 Y C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_1241_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X10 a_27_47# B2 a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VPWR B1 a_553_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 VGND A2 a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_553_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X14 a_27_47# B2 a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 VGND A2 a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 a_27_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 VGND A1 a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 Y C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X19 a_27_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 a_1241_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 VPWR B1 a_553_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X22 VPWR A1 a_1241_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 Y B2 a_553_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 a_1241_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X26 a_553_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 a_471_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X28 Y A2 a_1241_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 a_553_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X30 a_27_47# B1 a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X31 VGND A1 a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.11375 ps=1 w=0.65 l=0.15
X32 Y B2 a_553_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X33 a_1241_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X34 a_27_47# B1 a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X35 a_553_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X36 Y A2 a_1241_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X37 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X38 a_471_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X39 a_471_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21bai_1 VPWR VGND VPB VNB A1 B1_N Y A2
X0 a_388_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1275 pd=1.255 as=0.1525 ps=1.305 w=1 l=0.15
X1 a_105_352# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_297_47# a_105_352# Y VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_297_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 VPWR A1 a_388_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.1275 ps=1.255 w=1 l=0.15
X5 VGND A2 a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X6 VPWR B1_N a_105_352# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.17825 pd=1.4 as=0.1092 ps=1.36 w=0.42 l=0.15
X7 Y a_105_352# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.17825 ps=1.4 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a221oi_4 VPWR VGND VPB VNB C1 Y B2 B1 A2 A1
X0 Y A1 a_1241_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_453_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 Y B1 a_453_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25025 ps=1.42 w=0.65 l=0.15
X3 Y A1 a_1241_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 Y C1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 a_471_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.295 pd=2.59 as=0.135 ps=1.27 w=1 l=0.15
X6 Y B1 a_453_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VGND A2 a_1241_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_27_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR A2 a_471_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X11 a_453_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 a_471_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 VGND B2 a_453_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 a_1241_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 a_27_297# B2 a_471_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X16 a_453_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 a_1241_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 a_1241_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X21 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.09425 pd=0.94 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 VPWR A2 a_471_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 a_471_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X24 a_471_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 a_471_297# B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X26 VPWR A1 a_471_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 Y C1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X28 a_27_297# B1 a_471_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 VGND A2 a_1241_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X30 a_471_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X31 a_27_297# B1 a_471_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X32 a_1241_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.11375 ps=1 w=0.65 l=0.15
X33 a_471_297# B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X34 VPWR A1 a_471_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X35 a_27_297# B2 a_471_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X36 a_471_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X37 a_27_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X38 a_453_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.09425 ps=0.94 w=0.65 l=0.15
X39 VGND B2 a_453_47# VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor3_4 VGND VPWR VPB VNB B A Y C
X0 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_449_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_27_297# B a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 Y C a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_449_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 Y C a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X10 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_449_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X15 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 a_27_297# B a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 a_449_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X22 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X23 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor2_4 VGND VPWR VPB VNB Y B A
X0 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X6 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X11 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o41a_1 VGND VPWR VPB VNB X B1 A4 A3 A2 A1
X0 VGND A4 a_321_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_321_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.1235 ps=1.03 w=0.65 l=0.15
X2 a_103_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=1.52 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR a_103_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.425 ps=2.85 w=1 l=0.15
X4 VGND a_103_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.247 ps=2.06 w=0.65 l=0.15
X5 VGND A2 a_321_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X6 a_321_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.12675 ps=1.04 w=0.65 l=0.15
X7 a_511_297# A3 a_393_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.22 ps=1.44 w=1 l=0.15
X8 a_619_297# A2 a_511_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X9 a_321_47# B1 a_103_21# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10 a_393_297# A4 a_103_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.26 ps=1.52 w=1 l=0.15
X11 VPWR A1 a_619_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.195 ps=1.39 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfrtp_2 VGND VPWR VPB VNB CLK D RESET_B Q
X0 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X4 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X5 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X7 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X8 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X9 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X10 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X11 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X12 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X14 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X15 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X16 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X17 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X18 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X19 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X20 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X21 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X22 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X23 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X24 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X25 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X26 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X27 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X28 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X29 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
.ends

.subckt sky130_fd_sc_hd__and4bb_4 VGND VPWR VPB VNB A_N C D X B_N
X0 VPWR a_174_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X1 a_174_21# a_832_21# a_766_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X2 X a_174_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_832_21# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1764 ps=1.68 w=0.42 l=0.15
X4 a_766_47# a_27_47# a_652_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.1365 ps=1.07 w=0.65 l=0.15
X5 VPWR a_174_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 X a_174_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14075 ps=1.325 w=1 l=0.15
X7 VPWR B_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 a_652_47# C a_556_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1365 pd=1.07 as=0.10725 ps=0.98 w=0.65 l=0.15
X9 a_832_21# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.31165 ps=2.125 w=0.42 l=0.15
X10 X a_174_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X11 X a_174_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 a_556_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.11375 ps=1 w=0.65 l=0.15
X13 a_174_21# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.175 ps=1.35 w=1 l=0.15
X14 VPWR C a_174_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.165 ps=1.33 w=1 l=0.15
X15 VGND a_174_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 VGND a_174_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 VPWR a_832_21# a_174_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.31165 pd=2.125 as=0.165 ps=1.33 w=1 l=0.15
X18 a_174_21# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.21 ps=1.42 w=1 l=0.15
X19 VGND B_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__and4_4 VGND VPWR VPB VNB X D C B A
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_188_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.108875 pd=0.985 as=0.079625 ps=0.895 w=0.65 l=0.15
X3 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND D a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.141375 ps=1.085 w=0.65 l=0.15
X5 VPWR D a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.215 ps=1.43 w=1 l=0.15
X6 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X7 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.135 ps=1.27 w=1 l=0.15
X9 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.105625 ps=0.975 w=0.65 l=0.15
X10 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 a_27_47# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.215 pd=1.43 as=0.155 ps=1.31 w=1 l=0.15
X12 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X14 a_285_47# C a_188_47# VNB sky130_fd_pr__nfet_01v8 ad=0.141375 pd=1.085 as=0.108875 ps=0.985 w=0.65 l=0.15
X15 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.079625 pd=0.895 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o221ai_1 VGND VPWR VPB VNB A1 A2 Y B2 C1 B1
X0 a_109_47# B1 a_213_123# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1652 ps=1.82 w=0.65 l=0.15
X1 Y B2 a_295_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.12 ps=1.24 w=1 l=0.15
X2 VPWR A1 a_493_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3 a_213_123# B2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_295_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.12 pd=1.24 as=0.38 ps=1.76 w=1 l=0.15
X5 a_493_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.225 ps=1.45 w=1 l=0.15
X6 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.38 pd=1.76 as=0.28 ps=2.56 w=1 l=0.15
X7 VGND A2 a_213_123# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.117 ps=1.01 w=0.65 l=0.15
X8 a_213_123# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_109_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.1654 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a211oi_1 VPWR VGND VPB VNB Y C1 B1 A1 A2
X0 a_56_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VPWR A2 a_56_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
X3 a_139_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.2665 ps=2.12 w=0.65 l=0.15
X4 a_311_297# B1 a_56_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X5 Y C1 a_311_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X6 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X7 Y A1 a_139_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__dlxtn_2 VPWR VGND VPB VNB Q D GATE_N
X0 VPWR a_728_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 VGND a_728_21# a_663_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2 VPWR a_728_21# a_686_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VPWR GATE_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4 a_686_413# a_27_47# a_565_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.09555 ps=0.875 w=0.42 l=0.15
X5 VGND a_728_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 Q a_728_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1425 ps=1.285 w=1 l=0.15
X7 VGND a_565_413# a_728_21# VNB sky130_fd_pr__nfet_01v8 ad=0.092625 pd=0.935 as=0.169 ps=1.82 w=0.65 l=0.15
X8 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 a_663_47# a_193_47# a_565_413# VNB sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0504 ps=0.64 w=0.36 l=0.15
X10 a_469_369# a_303_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0968 pd=0.97 as=0.0864 ps=0.91 w=0.64 l=0.15
X11 VGND D a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X12 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X13 VPWR D a_303_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X14 a_565_413# a_193_47# a_469_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.09555 pd=0.875 as=0.0968 ps=0.97 w=0.42 l=0.15
X15 VPWR a_565_413# a_728_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1425 pd=1.285 as=0.26 ps=2.52 w=1 l=0.15
X16 a_469_47# a_303_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0777 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 VGND GATE_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X18 a_565_413# a_27_47# a_469_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0504 pd=0.64 as=0.0777 ps=0.81 w=0.36 l=0.15
X19 Q a_728_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.092625 ps=0.935 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand3_2 VGND VPWR VPB VNB C A Y B
X0 VGND C a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.2015 pd=1.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 a_277_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_27_47# B a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.31 pd=2.62 as=0.135 ps=1.27 w=1 l=0.15
X8 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 a_277_47# B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_8 VGND VPWR VPB VNB A X
X0 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X21 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o41ai_4 VGND VPWR VPB VNB B1 Y A4 A1 A2 A3
X0 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1 a_467_297# A4 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VPWR A1 a_1243_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 a_27_47# A4 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 Y A4 a_467_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 a_27_47# A4 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VGND A4 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 a_1243_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 VGND A4 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VPWR A1 a_1243_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X23 a_467_297# A4 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 a_1243_297# A2 a_885_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 Y A4 a_467_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X26 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X27 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X28 a_885_297# A2 a_1243_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X30 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X31 a_1243_297# A2 a_885_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X32 a_467_297# A3 a_885_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X33 a_885_297# A2 a_1243_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X34 a_885_297# A3 a_467_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X35 a_467_297# A3 a_885_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X36 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X37 a_1243_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X38 a_885_297# A3 a_467_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X39 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o211ai_2 VGND VPWR VPB VNB Y B1 A2 A1 C1
X0 a_286_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2 a_286_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.18525 ps=1.87 w=0.65 l=0.15
X3 Y A2 a_487_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4 VGND A1 a_286_47# VNB sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X5 Y C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.18525 ps=1.87 w=0.65 l=0.15
X6 VGND A2 a_286_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X7 a_487_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8 a_27_47# B1 a_286_47# VNB sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X9 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10 VPWR A1 a_487_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11 a_27_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X12 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X13 a_487_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X14 a_286_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X15 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__and4bb_1 VGND VPWR VPB VNB A_N B_N C D X
X0 VPWR D a_343_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.46 as=0.0777 ps=0.79 w=0.42 l=0.15
X1 a_223_47# B_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1386 pd=1.5 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 a_515_93# a_223_47# a_429_93# VNB sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 a_223_47# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1344 pd=1.48 as=0.0588 ps=0.7 w=0.42 l=0.15
X4 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.168 ps=1.64 w=0.42 l=0.15
X5 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.168 ps=1.64 w=0.42 l=0.15
X6 X a_343_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.172 ps=1.46 w=1 l=0.15
X7 a_429_93# a_27_47# a_343_93# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1176 ps=1.4 w=0.42 l=0.15
X8 VGND D a_615_93# VNB sky130_fd_pr__nfet_01v8 ad=0.1265 pd=1.11 as=0.0777 ps=0.79 w=0.42 l=0.15
X9 a_343_93# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X10 a_343_93# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X11 a_615_93# C a_515_93# VNB sky130_fd_pr__nfet_01v8 ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X12 X a_343_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1654 pd=1.82 as=0.1265 ps=1.11 w=0.65 l=0.15
X13 VPWR a_223_47# a_343_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand2_2 VGND VPWR VPB VNB Y A B
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3_4 VPWR VGND VPB VNB B C A X
X0 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.26 ps=1.45 w=0.65 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.4 ps=1.8 w=1 l=0.15
X2 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.20475 pd=1.93 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 VPWR A a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.4 pd=1.8 as=0.135 ps=1.27 w=1 l=0.15
X5 a_193_297# B a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.135 ps=1.27 w=1 l=0.15
X8 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 a_109_297# C a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13 VGND C a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o2111ai_1 VGND VPWR VPB VNB Y A1 A2 C1 D1 B1
X0 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.14 ps=1.28 w=1 l=0.15
X1 a_235_47# C1 a_163_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.06825 ps=0.86 w=0.65 l=0.15
X2 a_343_47# B1 a_235_47# VNB sky130_fd_pr__nfet_01v8 ad=0.131625 pd=1.055 as=0.12675 ps=1.04 w=0.65 l=0.15
X3 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2025 pd=1.405 as=0.195 ps=1.39 w=1 l=0.15
X4 a_454_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.2025 ps=1.405 w=1 l=0.15
X5 Y D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X6 VPWR A1 a_454_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.195 ps=1.39 w=1 l=0.15
X7 a_163_47# D1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X8 VGND A2 a_343_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.131625 ps=1.055 w=0.65 l=0.15
X9 a_343_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.12675 ps=1.04 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and3b_4 VGND VPWR VPB VNB A_N X B C
X0 a_98_199# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1491 pd=1.55 as=0.108375 ps=1.01 w=0.42 l=0.15
X1 X a_56_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2 VPWR a_56_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15825 pd=1.36 as=0.14 ps=1.28 w=1 l=0.15
X3 VGND a_56_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.108375 pd=1.01 as=0.091 ps=0.93 w=0.65 l=0.15
X4 VPWR a_98_199# a_56_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1875 pd=1.375 as=0.33 ps=2.66 w=1 l=0.15
X5 VPWR a_56_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.145 ps=1.29 w=1 l=0.15
X6 VGND a_56_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X7 a_257_47# B a_152_47# VNB sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.121875 ps=1.025 w=0.65 l=0.15
X8 X a_56_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X9 X a_56_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.1775 ps=1.355 w=1 l=0.15
X10 a_152_47# a_98_199# a_56_297# VNB sky130_fd_pr__nfet_01v8 ad=0.121875 pd=1.025 as=0.19825 ps=1.91 w=0.65 l=0.15
X11 VPWR C a_56_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.15 ps=1.3 w=1 l=0.15
X12 a_98_199# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1197 pd=1.41 as=0.15825 ps=1.36 w=0.42 l=0.15
X13 a_56_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.1875 ps=1.375 w=1 l=0.15
X14 VGND C a_257_47# VNB sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.07475 ps=0.88 w=0.65 l=0.15
X15 X a_56_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor3b_4 VGND VPWR VPB VNB A C_N B Y
X0 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 VPWR A a_197_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_555_297# a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 a_197_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VGND a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 a_197_297# B a_555_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8 VGND a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VGND C_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X12 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 Y a_27_47# a_555_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 Y a_27_47# a_555_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VPWR C_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X16 a_555_297# a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 a_555_297# B a_197_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 a_197_297# B a_555_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 a_555_297# B a_197_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X22 VPWR A a_197_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X23 a_197_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25675 ps=1.44 w=0.65 l=0.15
X25 Y a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a2111oi_4 VGND VPWR VPB VNB A1 Y D1 C1 A2 B1
X0 Y D1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1 a_455_297# B1 a_821_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.26 ps=2.52 w=1 l=0.15
X2 a_28_297# D1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 a_821_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X4 a_28_297# C1 a_455_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5 a_455_297# C1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 VGND D1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.091 ps=0.93 w=0.65 l=0.15
X7 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X8 VPWR A2 a_821_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.2 ps=1.4 w=1 l=0.15
X9 Y D1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X10 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X11 VGND D1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 Y D1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X13 a_821_297# B1 a_455_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X14 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X15 Y D1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X16 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.117 ps=1.01 w=0.65 l=0.15
X17 a_1205_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X18 a_28_297# C1 a_455_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14 ps=1.28 w=1 l=0.15
X19 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.12675 ps=1.04 w=0.65 l=0.15
X20 a_1205_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X21 a_821_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.14 ps=1.28 w=1 l=0.15
X22 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.091 ps=0.93 w=0.65 l=0.15
X23 Y A1 a_1205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X24 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X25 VPWR A1 a_821_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.145 ps=1.29 w=1 l=0.15
X26 Y A1 a_1205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.182 ps=1.86 w=0.65 l=0.15
X27 a_1205_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.121875 pd=1.025 as=0.091 ps=0.93 w=0.65 l=0.15
X28 a_28_297# D1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X29 VGND A2 a_1205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X30 a_455_297# B1 a_821_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X31 a_821_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2 pd=1.4 as=0.15 ps=1.3 w=1 l=0.15
X32 a_1205_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X33 VGND A2 a_1205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.121875 ps=1.025 w=0.65 l=0.15
X34 VPWR A1 a_821_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.14 ps=1.28 w=1 l=0.15
X35 a_821_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X36 VPWR A2 a_821_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X37 a_455_297# C1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X38 a_821_297# B1 a_455_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.14 ps=1.28 w=1 l=0.15
X39 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt dig_ctrl_top uio_in[4] clk ena rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4]
+ ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[5] uio_in[6]
+ uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6]
+ uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6]
+ uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6]
+ uo_out[7] clk_o port_ms_i port_ms_o[0] port_ms_o[1] port_ms_o[2] port_ms_o[3] port_ms_o[4]
+ port_ms_o[5] port_ms_o[6] port_ms_o[7] VDPWR VGND
X_2037_ VDPWR VGND VDPWR VGND _1010_ _0200_ _0741_ sky130_fd_sc_hd__and2_2
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[46\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[46\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[46\] clknet_leaf_16_clk sky130_fd_sc_hd__dlclkp_1
X_2106_ VDPWR VGND VDPWR VGND dig_ctrl_inst.cpu_inst.data\[4\] dig_ctrl_inst.cpu_inst.data\[6\]
+ dig_ctrl_inst.cpu_inst.data\[7\] dig_ctrl_inst.cpu_inst.data\[5\] _0799_ sky130_fd_sc_hd__or4_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[41\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[41\]\[3\] net221 dig_ctrl_inst.latch_mem_inst.gclk\[41\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_15_Left_93 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[30\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[30\]\[1\] net234 dig_ctrl_inst.latch_mem_inst.gclk\[30\]
+ sky130_fd_sc_hd__dlxtp_1
Xrebuffer7 VDPWR VGND VDPWR VGND net289 _1079_ sky130_fd_sc_hd__buf_2
X_1270_ VGND VDPWR VDPWR VGND _1118_ _1117_ _1114_ _1115_ _1116_ _1018_ sky130_fd_sc_hd__o41a_4
XFILLER_0_64_14 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
Xdig_ctrl_inst.latch_mem_inst.gen_words\[56\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[56\]\[6\] net196 dig_ctrl_inst.latch_mem_inst.gclk\[56\]
+ sky130_fd_sc_hd__dlxtp_1
X_1606_ VDPWR VGND VDPWR VGND _0315_ _0317_ _0316_ _0314_ _0318_ sky130_fd_sc_hd__or4_1
X_1468_ VDPWR VGND VDPWR VGND _0009_ _0194_ _0196_ sky130_fd_sc_hd__and2_1
Xfanout127 VGND VDPWR VDPWR VGND _1128_ net127 sky130_fd_sc_hd__clkbuf_2
Xfanout149 VDPWR VGND VDPWR VGND net149 net151 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout116 VDPWR VGND VDPWR VGND net117 net116 sky130_fd_sc_hd__buf_4
Xfanout105 VDPWR VGND VDPWR VGND _1134_ net105 sky130_fd_sc_hd__buf_4
Xfanout138 VDPWR VGND VDPWR VGND net138 _0227_ sky130_fd_sc_hd__buf_2
X_1537_ VGND VDPWR VDPWR VGND net171 net169 _0250_ sky130_fd_sc_hd__nor2_1
X_1399_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[57\] net148 _0154_
+ sky130_fd_sc_hd__and2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[45\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[45\]\[4\] net210 dig_ctrl_inst.latch_mem_inst.gclk\[45\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_64_125 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[34\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[34\]\[2\] net227 dig_ctrl_inst.latch_mem_inst.gclk\[34\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_0_Left_78 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_18_29 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[23\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[23\]\[0\] net247 dig_ctrl_inst.latch_mem_inst.gclk\[23\]
+ sky130_fd_sc_hd__dlxtp_1
X_2440_ VGND VDPWR VDPWR VGND clknet_leaf_6_clk _0048_ net145 dig_ctrl_inst.cpu_inst.r0\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_1253_ VGND VDPWR VDPWR VGND net257 _1101_ dig_ctrl_inst.cpu_inst.r1\[5\] sky130_fd_sc_hd__and2b_1
XFILLER_0_59_69 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1322_ VDPWR VGND VDPWR VGND _0119_ net129 net66 sky130_fd_sc_hd__and2_1
X_2371_ VDPWR VGND VDPWR VGND _0995_ net248 _0990_ _0111_ _0997_ sky130_fd_sc_hd__a22o_1
X_1184_ VDPWR VGND VDPWR VGND _1032_ dig_ctrl_inst.cpu_inst.r3\[3\] net256 net260
+ sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[11\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[11\]\[7\] net188 dig_ctrl_inst.latch_mem_inst.gclk\[11\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_46_136 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[5\].gen_latches\[0\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[5\]\[0\] net243 dig_ctrl_inst.latch_mem_inst.gclk\[5\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_27_Left_105 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[49\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[49\]\[5\] net199 dig_ctrl_inst.latch_mem_inst.gclk\[49\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_36_Left_114 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[38\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[38\]\[3\] net216 dig_ctrl_inst.latch_mem_inst.gclk\[38\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_45_Left_123 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[27\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[27\]\[1\] net237 dig_ctrl_inst.latch_mem_inst.gclk\[27\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_0_29 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_1871_ VGND VDPWR VDPWR VGND _0568_ _0287_ _0578_ _0577_ _0570_ sky130_fd_sc_hd__nor4_2
X_1940_ VDPWR VGND VDPWR VGND _0646_ net70 net74 dig_ctrl_inst.latch_mem_inst.RAM\[30\]\[6\]
+ sky130_fd_sc_hd__and3_2
XPHY_EDGE_ROW_54_Left_132 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_43_139 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_16_309 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_10_85 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2423_ VGND VDPWR VDPWR VGND clknet_leaf_13_clk _0031_ net139 dig_ctrl_inst.cpu_inst.instr\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_2354_ VGND VDPWR VDPWR VGND _0103_ net17 _0988_ dig_ctrl_inst.cpu_inst.port_o\[0\]
+ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_63_Left_141 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1236_ VGND VDPWR VDPWR VGND _1084_ _1083_ _1080_ _1081_ _1082_ _1018_ sky130_fd_sc_hd__o41a_4
X_2285_ VDPWR VGND VDPWR VGND _0830_ _0752_ _0833_ _0969_ sky130_fd_sc_hd__a21o_1
X_1305_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[9\] net150 _1143_
+ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_72_Left_150 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1167_ VGND VDPWR VDPWR VGND _1015_ net253 net252 dig_ctrl_inst.cpu_inst.instr\[6\]
+ dig_ctrl_inst.cpu_inst.instr\[7\] sky130_fd_sc_hd__or4b_4
XFILLER_0_19_169 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[9\].gen_latches\[1\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[9\]\[1\] net232 dig_ctrl_inst.latch_mem_inst.gclk\[9\]
+ sky130_fd_sc_hd__dlxtp_1
X_2070_ VGND VDPWR VDPWR VGND _0763_ _0762_ _1068_ _0761_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_3_Left_81 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1854_ VDPWR VGND VDPWR VGND _0129_ dig_ctrl_inst.latch_mem_inst.RAM\[13\]\[4\] _0114_
+ _0562_ dig_ctrl_inst.latch_mem_inst.RAM\[26\]\[4\] sky130_fd_sc_hd__a22o_1
X_1785_ VGND VDPWR VDPWR VGND _0135_ dig_ctrl_inst.latch_mem_inst.RAM\[33\]\[3\] _0491_
+ _0492_ _0493_ _0494_ sky130_fd_sc_hd__a2111o_1
X_1923_ VDPWR VGND VDPWR VGND _0629_ net112 net121 dig_ctrl_inst.latch_mem_inst.RAM\[2\]\[6\]
+ sky130_fd_sc_hd__and3_2
X_2406_ VGND VDPWR VDPWR VGND clknet_leaf_5_clk _0014_ net146 dig_ctrl_inst.cpu_inst.port_o\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_2337_ VGND VDPWR VDPWR VGND _0088_ net357 _0986_ dig_ctrl_inst.cpu_inst.port_o\[1\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_3 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
X_2268_ VGND VDPWR VDPWR VGND _0836_ _0908_ _0953_ _0954_ sky130_fd_sc_hd__o21a_1
X_2199_ VGND VDPWR VDPWR VGND _0887_ _0770_ _0837_ _0836_ _0888_ _0886_ sky130_fd_sc_hd__o221a_1
X_1219_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.r0\[0\] _1019_ _1066_ _1065_
+ _1067_ sky130_fd_sc_hd__o22a_2
XFILLER_0_22_109 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[53\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[53\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[53\] clknet_leaf_17_clk sky130_fd_sc_hd__dlclkp_1
Xhold52 VGND VDPWR VDPWR VGND net334 dig_ctrl_inst.synchronizer_port_i_inst\[2\].pipe\[0\]
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 VGND VDPWR VDPWR VGND net356 dig_ctrl_inst.spi_data_i\[5\] sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 VGND VDPWR VDPWR VGND net345 dig_ctrl_inst.spi_receiver_inst.spi_mosi_sync
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 VGND VDPWR VDPWR VGND net323 dig_ctrl_inst.latch_mem_inst.wdata\[4\] sky130_fd_sc_hd__dlygate4sd3_1
Xhold96 VGND VDPWR VDPWR VGND net378 dig_ctrl_inst.cpu_inst.r2\[4\] sky130_fd_sc_hd__dlygate4sd3_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[60\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[60\]\[1\] net234 dig_ctrl_inst.latch_mem_inst.gclk\[60\]
+ sky130_fd_sc_hd__dlxtp_1
Xhold85 VGND VDPWR VDPWR VGND net367 dig_ctrl_inst.cpu_inst.r1\[1\] sky130_fd_sc_hd__dlygate4sd3_1
X_1570_ VGND VDPWR VDPWR VGND _0282_ net82 net119 net123 net68 net130 sky130_fd_sc_hd__a32o_1
XANTENNA_5 VGND VDPWR VDPWR VGND _0560_ sky130_fd_sc_hd__diode_2
XFILLER_0_21_164 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xrebuffer17 VDPWR VGND VDPWR VGND net299 net300 sky130_fd_sc_hd__dlygate4sd1_1
X_2122_ VDPWR VGND VDPWR VGND _0814_ net137 net138 net157 sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[52\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[52\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[52\] sky130_fd_sc_hd__clkbuf_4
X_2053_ VGND VDPWR VDPWR VGND _0746_ net254 _1015_ _0744_ _0745_ sky130_fd_sc_hd__o211a_1
X_2528__275 VGND VDPWR VDPWR VGND net275 _2528__275/HI sky130_fd_sc_hd__conb_1
X_1837_ VGND VDPWR VDPWR VGND _0545_ net58 net92 net108 dig_ctrl_inst.latch_mem_inst.RAM\[43\]\[4\]
+ sky130_fd_sc_hd__and4_1
X_1906_ VDPWR VGND VDPWR VGND _0613_ net52 net76 dig_ctrl_inst.latch_mem_inst.RAM\[44\]\[5\]
+ sky130_fd_sc_hd__and3_2
X_1768_ VGND VDPWR VDPWR VGND _0153_ dig_ctrl_inst.latch_mem_inst.RAM\[55\]\[3\] _0474_
+ _0475_ _0476_ _0477_ sky130_fd_sc_hd__a2111o_1
X_1699_ VDPWR VGND VDPWR VGND _0409_ net85 net126 dig_ctrl_inst.latch_mem_inst.RAM\[10\]\[2\]
+ sky130_fd_sc_hd__and3_2
XFILLER_0_12_197 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xoutput20 VDPWR VGND VDPWR VGND port_ms_o[3] net20 sky130_fd_sc_hd__buf_2
Xoutput31 VDPWR VGND VDPWR VGND uo_out[3] net31 sky130_fd_sc_hd__buf_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[53\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[53\]\[0\] net242 dig_ctrl_inst.latch_mem_inst.gclk\[53\]
+ sky130_fd_sc_hd__dlxtp_1
X_1622_ VGND VDPWR VDPWR VGND _1143_ dig_ctrl_inst.latch_mem_inst.RAM\[9\]\[0\] _0295_
+ _0299_ _0304_ _0334_ sky130_fd_sc_hd__a2111o_1
X_1553_ VGND VDPWR VDPWR VGND _0266_ _0252_ net167 net166 sky130_fd_sc_hd__nand3b_1
X_1484_ VDPWR VGND VDPWR VGND _0173_ dig_ctrl_inst.cpu_inst.skip _0202_ _0203_ sky130_fd_sc_hd__a21o_1
X_2105_ VGND VDPWR VDPWR VGND _0798_ _0797_ _0796_ _0789_ _0782_ sky130_fd_sc_hd__and4_1
X_2036_ VGND VDPWR VDPWR VGND _0033_ _0740_ _0276_ dig_ctrl_inst.cpu_inst.instr\[7\]
+ sky130_fd_sc_hd__mux2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[41\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[41\]\[7\] net184 dig_ctrl_inst.latch_mem_inst.gclk\[41\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[30\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[30\]\[5\] net205 dig_ctrl_inst.latch_mem_inst.gclk\[30\]
+ sky130_fd_sc_hd__dlxtp_1
Xrebuffer8 VDPWR VGND VDPWR VGND net290 net291 sky130_fd_sc_hd__dlymetal6s4s_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[57\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[57\]\[1\] net232 dig_ctrl_inst.latch_mem_inst.gclk\[57\]
+ sky130_fd_sc_hd__dlxtp_1
X_1605_ VDPWR VGND VDPWR VGND _0137_ dig_ctrl_inst.latch_mem_inst.RAM\[16\]\[0\] _0119_
+ _0317_ dig_ctrl_inst.latch_mem_inst.RAM\[35\]\[0\] sky130_fd_sc_hd__a22o_1
X_1536_ VGND VDPWR VDPWR VGND net170 _0249_ net169 sky130_fd_sc_hd__nand2_1
Xfanout117 VDPWR VGND VDPWR VGND _1129_ net117 sky130_fd_sc_hd__buf_4
XFILLER_0_38_60 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
Xfanout106 VDPWR VGND VDPWR VGND net107 net106 sky130_fd_sc_hd__buf_4
X_1467_ VGND VDPWR VDPWR VGND _1096_ _0195_ _0184_ _0196_ sky130_fd_sc_hd__o21a_1
Xfanout128 VGND VDPWR VDPWR VGND net130 net128 sky130_fd_sc_hd__clkbuf_2
Xfanout139 VGND VDPWR VDPWR VGND net140 net139 sky130_fd_sc_hd__clkbuf_4
X_1398_ VGND VDPWR VDPWR VGND _0154_ net114 net90 net42 sky130_fd_sc_hd__and3_4
X_2019_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[3\]\[7\] _1135_ _0724_
+ _0120_ dig_ctrl_inst.latch_mem_inst.RAM\[17\]\[7\] _0723_ sky130_fd_sc_hd__a221o_1
XFILLER_0_54_81 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[1\].gen_latches\[3\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[1\]\[3\] net220 dig_ctrl_inst.latch_mem_inst.gclk\[1\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[34\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[34\]\[6\] net191 dig_ctrl_inst.latch_mem_inst.gclk\[34\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[23\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[23\]\[4\] net211 dig_ctrl_inst.latch_mem_inst.gclk\[23\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_50_17 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_59_48 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_2370_ VGND VDPWR VDPWR VGND _0990_ _0996_ _0997_ sky130_fd_sc_hd__nor2_1
X_1321_ VGND VDPWR VDPWR VGND _1112_ _0118_ _1127_ sky130_fd_sc_hd__and2b_1
X_1252_ VDPWR VGND VDPWR VGND _1100_ dig_ctrl_inst.cpu_inst.r3\[5\] net257 net261
+ sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[12\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[12\]\[2\] net231 dig_ctrl_inst.latch_mem_inst.gclk\[12\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[45\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[45\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[45\] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_73 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1183_ VGND VDPWR VDPWR VGND net258 _1031_ net254 sky130_fd_sc_hd__nand2_1
X_2499_ VGND VDPWR VDPWR VGND clknet_leaf_5_clk _0096_ net177 net29 sky130_fd_sc_hd__dfrtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[58\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[58\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[58\] clknet_leaf_1_clk sky130_fd_sc_hd__dlclkp_1
XFILLER_0_64_3 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_12_Right_12 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1519_ VDPWR VGND VDPWR VGND _0998_ dig_ctrl_inst.cpu_inst.r2\[7\] _0232_ dig_ctrl_inst.cpu_inst.r1\[7\]
+ _1022_ net299 sky130_fd_sc_hd__a221o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[5\].gen_latches\[4\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[5\]\[4\] net213 dig_ctrl_inst.latch_mem_inst.gclk\[5\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_21_Right_21 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_37_148 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_181 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_Right_30 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[38\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[38\]\[7\] net184 dig_ctrl_inst.latch_mem_inst.gclk\[38\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[27\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[27\]\[5\] net204 dig_ctrl_inst.latch_mem_inst.gclk\[27\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[60\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[60\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[60\] clknet_leaf_0_clk sky130_fd_sc_hd__dlclkp_1
X_1870_ VDPWR VGND VDPWR VGND _0575_ _0576_ _0574_ _0577_ sky130_fd_sc_hd__or3_1
XFILLER_0_36_181 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_2353_ VDPWR VGND VDPWR VGND _0800_ _0988_ dig_ctrl_inst.cpu_inst.data\[0\] dig_ctrl_inst.cpu_inst.port_stb_o
+ _0801_ sky130_fd_sc_hd__nand4_4
X_2422_ VGND VDPWR VDPWR VGND clknet_leaf_13_clk _0030_ net139 dig_ctrl_inst.cpu_inst.instr\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[16\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[16\]\[3\] net217 dig_ctrl_inst.latch_mem_inst.gclk\[16\]
+ sky130_fd_sc_hd__dlxtp_1
X_1166_ VGND VDPWR VDPWR VGND net252 net253 _1014_ sky130_fd_sc_hd__nand2b_1
X_2284_ VGND VDPWR VDPWR VGND _0053_ _0968_ _0967_ net374 sky130_fd_sc_hd__mux2_1
X_1235_ VDPWR VGND VDPWR VGND net255 dig_ctrl_inst.cpu_inst.r0\[1\] net259 _1083_
+ sky130_fd_sc_hd__or3_1
X_1304_ VGND VDPWR VDPWR VGND _1143_ net120 net116 net90 sky130_fd_sc_hd__and3_4
X_1999_ VDPWR VGND VDPWR VGND _0704_ net43 net129 dig_ctrl_inst.latch_mem_inst.RAM\[48\]\[7\]
+ sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[9\].gen_latches\[5\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[9\]\[5\] net200 dig_ctrl_inst.latch_mem_inst.gclk\[9\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[2\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[2\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[2\] sky130_fd_sc_hd__clkbuf_4
X_1922_ VDPWR VGND VDPWR VGND _0628_ net43 net129 dig_ctrl_inst.latch_mem_inst.RAM\[48\]\[6\]
+ sky130_fd_sc_hd__and3_2
X_1784_ VGND VDPWR VDPWR VGND _0493_ net62 net99 net103 dig_ctrl_inst.latch_mem_inst.RAM\[23\]\[3\]
+ sky130_fd_sc_hd__and4_1
X_1853_ VDPWR VGND VDPWR VGND _0135_ dig_ctrl_inst.latch_mem_inst.RAM\[21\]\[4\] _0124_
+ _0561_ dig_ctrl_inst.latch_mem_inst.RAM\[33\]\[4\] sky130_fd_sc_hd__a22o_1
X_2336_ VGND VDPWR VDPWR VGND _0087_ net380 _0986_ dig_ctrl_inst.cpu_inst.port_o\[0\]
+ sky130_fd_sc_hd__mux2_1
X_2405_ VGND VDPWR VDPWR VGND clknet_leaf_6_clk _0013_ net146 dig_ctrl_inst.cpu_inst.port_o\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_2267_ VGND VDPWR VDPWR VGND _0952_ _0770_ _0817_ _0768_ _0953_ _0886_ sky130_fd_sc_hd__o221a_1
X_2198_ VGND VDPWR VDPWR VGND _0887_ _0776_ _1068_ _0761_ sky130_fd_sc_hd__mux2_1
X_1218_ VGND VDPWR VDPWR VGND net258 _1066_ dig_ctrl_inst.cpu_inst.r2\[0\] sky130_fd_sc_hd__and2b_1
X_1149_ VDPWR VGND VDPWR VGND _0998_ net265 sky130_fd_sc_hd__inv_2
XFILLER_0_30_165 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xhold86 VGND VDPWR VDPWR VGND net368 dig_ctrl_inst.cpu_inst.r3\[5\] sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 VGND VDPWR VDPWR VGND net357 dig_ctrl_inst.spi_data_i\[1\] sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 VGND VDPWR VDPWR VGND net324 dig_ctrl_inst.latch_mem_inst.wdata\[2\] sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 VGND VDPWR VDPWR VGND net346 dig_ctrl_inst.cpu_inst.prev_state\[0\] sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 VGND VDPWR VDPWR VGND net335 dig_ctrl_inst.synchronizer_mode_i_inst.pipe\[0\]
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 VGND VDPWR VDPWR VGND net379 dig_ctrl_inst.cpu_inst.r2\[0\] sky130_fd_sc_hd__dlygate4sd3_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[60\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[60\]\[5\] net203 dig_ctrl_inst.latch_mem_inst.gclk\[60\]
+ sky130_fd_sc_hd__dlxtp_1
XANTENNA_6 VGND VDPWR VDPWR VGND _0592_ sky130_fd_sc_hd__diode_2
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[38\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[38\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[38\] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_21_154 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_16_41 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2052_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.instr\[7\] dig_ctrl_inst.cpu_inst.instr\[6\]
+ _0745_ sky130_fd_sc_hd__nand2b_1
X_2121_ VDPWR VGND VDPWR VGND _0813_ _0812_ _0810_ _0772_ sky130_fd_sc_hd__and3_2
XFILLER_0_76_338 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_32_95 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1905_ VDPWR VGND VDPWR VGND _0612_ net61 net93 dig_ctrl_inst.latch_mem_inst.RAM\[22\]\[5\]
+ sky130_fd_sc_hd__and3_2
X_1836_ VDPWR VGND VDPWR VGND _0544_ net72 net123 dig_ctrl_inst.latch_mem_inst.RAM\[14\]\[4\]
+ sky130_fd_sc_hd__and3_2
XPHY_EDGE_ROW_6_Right_6 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1698_ VDPWR VGND VDPWR VGND _0408_ net87 net122 dig_ctrl_inst.latch_mem_inst.RAM\[8\]\[2\]
+ sky130_fd_sc_hd__and3_2
X_1767_ VGND VDPWR VDPWR VGND _0476_ net51 net102 net131 dig_ctrl_inst.latch_mem_inst.RAM\[35\]\[3\]
+ sky130_fd_sc_hd__and4_1
X_2319_ VGND VDPWR VDPWR VGND _0980_ dig_ctrl_inst.spi_data_i\[2\] dig_ctrl_inst.spi_receiver_inst.spi_cnt\[0\]
+ dig_ctrl_inst.spi_data_i\[3\] sky130_fd_sc_hd__mux2_1
Xoutput21 VDPWR VGND VDPWR VGND port_ms_o[4] net21 sky130_fd_sc_hd__buf_2
Xoutput32 VDPWR VGND VDPWR VGND uo_out[4] net32 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_59_Right_59 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1621_ VGND VDPWR VDPWR VGND _0141_ dig_ctrl_inst.latch_mem_inst.RAM\[41\]\[0\] _0292_
+ _0298_ _0303_ _0333_ sky130_fd_sc_hd__a2111o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[53\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[53\]\[4\] net208 dig_ctrl_inst.latch_mem_inst.gclk\[53\]
+ sky130_fd_sc_hd__dlxtp_1
X_1552_ VDPWR VGND VDPWR VGND _0264_ _0257_ _0263_ _0265_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_68_Right_68 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2104_ VGND VDPWR VDPWR VGND _0793_ _0258_ _0785_ _0259_ _0797_ _0795_ sky130_fd_sc_hd__o221a_1
X_1483_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.cpu_state\[1\] _0999_ _0202_
+ net248 sky130_fd_sc_hd__o21ai_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[42\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[42\]\[2\] net230 dig_ctrl_inst.latch_mem_inst.gclk\[42\]
+ sky130_fd_sc_hd__dlxtp_1
X_2035_ VGND VDPWR VDPWR VGND _0740_ _0728_ _0739_ _0729_ _0686_ sky130_fd_sc_hd__o31a_1
XPHY_EDGE_ROW_77_Right_77 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_17_213 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
Xdig_ctrl_inst.latch_mem_inst.gen_words\[31\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[31\]\[0\] net246 dig_ctrl_inst.latch_mem_inst.gclk\[31\]
+ sky130_fd_sc_hd__dlxtp_1
X_1819_ VGND VDPWR VDPWR VGND _0151_ dig_ctrl_inst.latch_mem_inst.RAM\[53\]\[4\] _0524_
+ _0525_ _0526_ _0527_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_4_162 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_7_50 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_67_113 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xrebuffer9 VGND VDPWR VDPWR VGND net291 net302 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_290 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_17 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_3_19 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[57\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[57\]\[5\] net202 dig_ctrl_inst.latch_mem_inst.gclk\[57\]
+ sky130_fd_sc_hd__dlxtp_1
Xfanout107 VDPWR VGND VDPWR VGND net108 net107 sky130_fd_sc_hd__buf_4
X_1604_ VGND VDPWR VDPWR VGND _0316_ net59 net98 dig_ctrl_inst.latch_mem_inst.RAM\[36\]\[0\]
+ _0114_ dig_ctrl_inst.latch_mem_inst.RAM\[13\]\[0\] sky130_fd_sc_hd__a32o_1
Xfanout118 VGND VDPWR VDPWR VGND net119 net118 sky130_fd_sc_hd__clkbuf_2
X_1535_ VGND VDPWR VDPWR VGND _0246_ _0248_ _0247_ sky130_fd_sc_hd__nand2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[46\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[46\]\[3\] net217 dig_ctrl_inst.latch_mem_inst.gclk\[46\]
+ sky130_fd_sc_hd__dlxtp_1
Xfanout129 VGND VDPWR VDPWR VGND net130 net129 sky130_fd_sc_hd__clkbuf_2
X_1466_ VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_addr\[3\] dig_ctrl_inst.spi_addr\[4\]
+ _0195_ _0191_ sky130_fd_sc_hd__nand3_1
X_1397_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[56\] net48 net88
+ net153 sky130_fd_sc_hd__and3_2
X_2018_ VDPWR VGND VDPWR VGND _0279_ dig_ctrl_inst.latch_mem_inst.RAM\[32\]\[7\] _0134_
+ _0723_ dig_ctrl_inst.latch_mem_inst.RAM\[6\]\[7\] sky130_fd_sc_hd__a22o_1
XFILLER_0_54_93 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[35\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[35\]\[1\] net235 dig_ctrl_inst.latch_mem_inst.gclk\[35\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[1\].gen_latches\[7\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[1\]\[7\] net185 dig_ctrl_inst.latch_mem_inst.gclk\[1\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_13_260 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_1320_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[15\] net155 _0117_
+ sky130_fd_sc_hd__and2_1
X_1182_ VGND VDPWR VDPWR VGND _1025_ _1030_ _1010_ sky130_fd_sc_hd__and2_4
X_1251_ VGND VDPWR VDPWR VGND net257 net260 _1099_ dig_ctrl_inst.cpu_inst.r2\[5\]
+ sky130_fd_sc_hd__and3b_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[12\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[12\]\[6\] net191 dig_ctrl_inst.latch_mem_inst.gclk\[12\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_24_85 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_40_73 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2498_ VGND VDPWR VDPWR VGND clknet_leaf_5_clk _0095_ net177 net28 sky130_fd_sc_hd__dfrtp_1
X_1449_ VGND VDPWR VDPWR VGND _0182_ _0183_ _0003_ sky130_fd_sc_hd__nor2_1
XFILLER_0_57_3 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1518_ VDPWR VGND VDPWR VGND _0231_ dig_ctrl_inst.cpu_inst.r3\[7\] net262 net265
+ sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[39\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[39\]\[2\] net231 dig_ctrl_inst.latch_mem_inst.gclk\[39\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_5_290 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[28\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[28\]\[0\] net240 dig_ctrl_inst.latch_mem_inst.gclk\[28\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_36_193 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1303_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[8\] net89 net126
+ net155 sky130_fd_sc_hd__and3_2
X_2352_ VGND VDPWR VDPWR VGND _0102_ net35 _0987_ dig_ctrl_inst.cpu_inst.port_o\[7\]
+ sky130_fd_sc_hd__mux2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[16\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[16\]\[7\] net184 dig_ctrl_inst.latch_mem_inst.gclk\[16\]
+ sky130_fd_sc_hd__dlxtp_1
X_2283_ VGND VDPWR VDPWR VGND _0751_ _0798_ _0968_ net164 sky130_fd_sc_hd__o21ai_1
X_2421_ VGND VDPWR VDPWR VGND clknet_leaf_9_clk _0029_ net141 dig_ctrl_inst.cpu_inst.arg1\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_40 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1165_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.instr\[6\] dig_ctrl_inst.cpu_inst.instr\[7\]
+ _1013_ sky130_fd_sc_hd__nor2_1
X_1234_ VGND VDPWR VDPWR VGND net255 _1082_ dig_ctrl_inst.cpu_inst.r1\[1\] sky130_fd_sc_hd__and2b_1
XFILLER_0_27_160 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_1998_ VDPWR VGND VDPWR VGND _0703_ net70 net83 dig_ctrl_inst.latch_mem_inst.RAM\[26\]\[7\]
+ sky130_fd_sc_hd__and3_2
XFILLER_0_42_141 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xwire113 VGND VDPWR VDPWR VGND net113 _1132_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_119 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
X_1852_ VDPWR VGND VDPWR VGND _0159_ dig_ctrl_inst.latch_mem_inst.RAM\[15\]\[4\] _0117_
+ _0560_ dig_ctrl_inst.latch_mem_inst.RAM\[62\]\[4\] sky130_fd_sc_hd__a22o_1
X_1921_ VGND VDPWR VDPWR VGND _0627_ net66 net104 net133 dig_ctrl_inst.latch_mem_inst.RAM\[19\]\[6\]
+ sky130_fd_sc_hd__and4_1
XFILLER_0_16_108 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1783_ VDPWR VGND VDPWR VGND _0492_ net110 net122 dig_ctrl_inst.latch_mem_inst.RAM\[2\]\[3\]
+ sky130_fd_sc_hd__and3_2
X_2404_ VGND VDPWR VDPWR VGND clknet_leaf_6_clk _0012_ net146 dig_ctrl_inst.cpu_inst.port_o\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_2335_ VGND VDPWR VDPWR VGND _0804_ _0986_ dig_ctrl_inst.cpu_inst.port_stb_o sky130_fd_sc_hd__nand2_4
X_2266_ VGND VDPWR VDPWR VGND _0814_ _0952_ _0817_ sky130_fd_sc_hd__and2b_1
X_2197_ VGND VDPWR VDPWR VGND net168 _0886_ _0769_ sky130_fd_sc_hd__nand2_1
X_1217_ VGND VDPWR VDPWR VGND _1065_ _1064_ _1000_ dig_ctrl_inst.cpu_inst.r1\[0\]
+ _1018_ sky130_fd_sc_hd__a211o_1
XFILLER_0_15_163 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[61\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[61\]\[0\] net242 dig_ctrl_inst.latch_mem_inst.gclk\[61\]
+ sky130_fd_sc_hd__dlxtp_1
Xhold98 VGND VDPWR VDPWR VGND net380 dig_ctrl_inst.spi_data_i\[0\] sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 VGND VDPWR VDPWR VGND net336 dig_ctrl_inst.spi_receiver_inst.synchronizer_spi_mosi.pipe\[0\]
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 VGND VDPWR VDPWR VGND net347 _0042_ sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 VGND VDPWR VDPWR VGND net325 dig_ctrl_inst.latch_mem_inst.wdata\[0\] sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 VGND VDPWR VDPWR VGND net369 dig_ctrl_inst.cpu_inst.r1\[2\] sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 VGND VDPWR VDPWR VGND net358 dig_ctrl_inst.cpu_inst.r3\[1\] sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_7 VGND VDPWR VDPWR VGND _0666_ sky130_fd_sc_hd__diode_2
X_2120_ VGND VDPWR VDPWR VGND _0768_ _0808_ _0765_ _0811_ _0812_ sky130_fd_sc_hd__o22a_1
Xrebuffer19 VDPWR VGND VDPWR VGND net301 _1094_ sky130_fd_sc_hd__dlygate4sd1_1
X_2051_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.instr\[6\] _0744_ dig_ctrl_inst.cpu_inst.instr\[7\]
+ sky130_fd_sc_hd__nand2b_2
X_1835_ VDPWR VGND VDPWR VGND _0543_ net58 net95 dig_ctrl_inst.latch_mem_inst.RAM\[38\]\[4\]
+ sky130_fd_sc_hd__and3_2
X_1904_ VGND VDPWR VDPWR VGND _0117_ dig_ctrl_inst.latch_mem_inst.RAM\[15\]\[5\] _0608_
+ _0609_ _0610_ _0611_ sky130_fd_sc_hd__a2111o_1
X_1697_ VDPWR VGND VDPWR VGND _0407_ net71 net97 dig_ctrl_inst.latch_mem_inst.RAM\[20\]\[2\]
+ sky130_fd_sc_hd__and3_2
X_1766_ VDPWR VGND VDPWR VGND _0475_ net53 net93 dig_ctrl_inst.latch_mem_inst.RAM\[38\]\[3\]
+ sky130_fd_sc_hd__and3_2
X_2318_ VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_data_i\[6\] dig_ctrl_inst.spi_data_i\[7\]
+ dig_ctrl_inst.spi_receiver_inst.spi_cnt\[0\] dig_ctrl_inst.spi_data_i\[4\] dig_ctrl_inst.spi_data_i\[5\]
+ dig_ctrl_inst.spi_receiver_inst.spi_cnt\[1\] _0979_ sky130_fd_sc_hd__mux4_1
X_2249_ VGND VDPWR VDPWR VGND _0936_ _0749_ _0935_ _0747_ sky130_fd_sc_hd__mux2_1
Xoutput22 VDPWR VGND VDPWR VGND port_ms_o[5] net22 sky130_fd_sc_hd__buf_2
Xoutput33 VDPWR VGND VDPWR VGND uo_out[5] net33 sky130_fd_sc_hd__buf_2
XFILLER_0_9_3 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_41_206 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1482_ VGND VDPWR VDPWR VGND _0200_ _1027_ _0201_ sky130_fd_sc_hd__nand2b_1
X_1551_ VGND VDPWR VDPWR VGND _1068_ _0264_ net164 sky130_fd_sc_hd__nand2_1
X_1620_ VGND VDPWR VDPWR VGND _0135_ dig_ctrl_inst.latch_mem_inst.RAM\[33\]\[0\] _0291_
+ _0296_ _0297_ _0332_ sky130_fd_sc_hd__a2111o_1
X_2103_ VGND VDPWR VDPWR VGND _0796_ net164 _0750_ _0784_ _0794_ sky130_fd_sc_hd__o211a_1
X_2034_ VDPWR VGND VDPWR VGND _0738_ _0734_ _0719_ _0287_ _0739_ sky130_fd_sc_hd__or4_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[42\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[42\]\[6\] net198 dig_ctrl_inst.latch_mem_inst.gclk\[42\]
+ sky130_fd_sc_hd__dlxtp_1
X_1818_ VDPWR VGND VDPWR VGND _0526_ net54 net96 dig_ctrl_inst.latch_mem_inst.RAM\[36\]\[4\]
+ sky130_fd_sc_hd__and3_2
X_1749_ VDPWR VGND VDPWR VGND _0455_ _0457_ _0456_ _0454_ _0458_ sky130_fd_sc_hd__or4_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[31\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[31\]\[4\] net208 dig_ctrl_inst.latch_mem_inst.gclk\[31\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_63_331 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[20\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[20\]\[2\] net228 dig_ctrl_inst.latch_mem_inst.gclk\[20\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_48_29 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
Xdig_ctrl_inst.latch_mem_inst.gen_words\[58\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[58\]\[0\] net246 dig_ctrl_inst.latch_mem_inst.gclk\[58\]
+ sky130_fd_sc_hd__dlxtp_1
Xfanout119 VGND VDPWR VDPWR VGND _1129_ net119 sky130_fd_sc_hd__clkbuf_4
X_1465_ VGND VDPWR VDPWR VGND _0194_ _0191_ _0185_ dig_ctrl_inst.spi_addr\[3\] dig_ctrl_inst.spi_addr\[4\]
+ sky130_fd_sc_hd__a31o_1
Xfanout108 VDPWR VGND VDPWR VGND _1134_ net108 sky130_fd_sc_hd__buf_4
X_1603_ VDPWR VGND VDPWR VGND _0155_ dig_ctrl_inst.latch_mem_inst.RAM\[21\]\[0\] _0124_
+ _0315_ dig_ctrl_inst.latch_mem_inst.RAM\[58\]\[0\] sky130_fd_sc_hd__a22o_1
X_1534_ VGND VDPWR VDPWR VGND _0247_ net167 net166 sky130_fd_sc_hd__or2_1
X_2017_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[25\]\[7\] _0128_ _0722_
+ _0139_ dig_ctrl_inst.latch_mem_inst.RAM\[39\]\[7\] _0721_ sky130_fd_sc_hd__a221o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[2\].gen_latches\[2\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[2\]\[2\] net225 dig_ctrl_inst.latch_mem_inst.gclk\[2\]
+ sky130_fd_sc_hd__dlxtp_1
X_1396_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[55\] net149 _0153_
+ sky130_fd_sc_hd__and2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[46\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[46\]\[7\] net183 dig_ctrl_inst.latch_mem_inst.gclk\[46\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_64_106 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_19_Left_97 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_13_272 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
Xdig_ctrl_inst.latch_mem_inst.gen_words\[35\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[35\]\[5\] net200 dig_ctrl_inst.latch_mem_inst.gclk\[35\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[24\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[24\]\[3\] net216 dig_ctrl_inst.latch_mem_inst.gclk\[24\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[11\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[11\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[11\] clknet_leaf_1_clk sky130_fd_sc_hd__dlclkp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[13\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[13\]\[1\] net236 dig_ctrl_inst.latch_mem_inst.gclk\[13\]
+ sky130_fd_sc_hd__dlxtp_1
X_1181_ VGND VDPWR VDPWR VGND _1029_ dig_ctrl_inst.cpu_inst.ip\[3\] _1027_ net292
+ net182 sky130_fd_sc_hd__o211a_4
X_1250_ VGND VDPWR VDPWR VGND _1098_ net182 net297 _1027_ dig_ctrl_inst.cpu_inst.ip\[5\]
+ sky130_fd_sc_hd__o211a_1
X_1448_ VDPWR VGND VDPWR VGND _0181_ dig_ctrl_inst.spi_receiver_inst.spi_cnt\[0\]
+ dig_ctrl_inst.spi_receiver_inst.spi_cnt\[1\] _0183_ sky130_fd_sc_hd__a21oi_1
X_2497_ VGND VDPWR VDPWR VGND clknet_leaf_8_clk dig_ctrl_inst.cpu_inst.stb_o net180
+ dig_ctrl_inst.stb_d sky130_fd_sc_hd__dfrtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[6\].gen_latches\[3\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[6\]\[3\] net220 dig_ctrl_inst.latch_mem_inst.gclk\[6\]
+ sky130_fd_sc_hd__dlxtp_1
X_1517_ VGND VDPWR VDPWR VGND _0230_ _0228_ _0229_ sky130_fd_sc_hd__or2_1
X_1379_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[46\] net51 net72
+ net148 sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[39\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[39\]\[6\] net191 dig_ctrl_inst.latch_mem_inst.gclk\[39\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[28\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[28\]\[4\] net209 dig_ctrl_inst.latch_mem_inst.gclk\[28\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[17\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[17\]\[2\] net230 dig_ctrl_inst.latch_mem_inst.gclk\[17\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_43_109 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xfanout90 VGND VDPWR VDPWR VGND net92 net90 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_23_Left_101 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2420_ VGND VDPWR VDPWR VGND clknet_leaf_9_clk _0028_ net141 dig_ctrl_inst.cpu_inst.arg1\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_2351_ VGND VDPWR VDPWR VGND _0101_ net34 _0987_ dig_ctrl_inst.cpu_inst.port_o\[6\]
+ sky130_fd_sc_hd__mux2_1
X_1302_ VDPWR VGND VDPWR VGND net124 net88 _1142_ sky130_fd_sc_hd__and2_2
X_1233_ VGND VDPWR VDPWR VGND net255 net259 _1081_ dig_ctrl_inst.cpu_inst.r2\[1\]
+ sky130_fd_sc_hd__and3b_1
X_2282_ VGND VDPWR VDPWR VGND _0967_ _1022_ _0175_ _0756_ sky130_fd_sc_hd__and3_4
XPHY_EDGE_ROW_32_Left_110 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1164_ VDPWR VGND VDPWR VGND _1012_ _1011_ sky130_fd_sc_hd__inv_2
X_1997_ VDPWR VGND VDPWR VGND _0702_ net49 net85 dig_ctrl_inst.latch_mem_inst.RAM\[58\]\[7\]
+ sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[41\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[41\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[41\] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_21_337 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1851_ VDPWR VGND VDPWR VGND _0152_ dig_ctrl_inst.latch_mem_inst.RAM\[47\]\[4\] _0146_
+ _0559_ dig_ctrl_inst.latch_mem_inst.RAM\[54\]\[4\] sky130_fd_sc_hd__a22o_1
XFILLER_0_8_309 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
X_1920_ VGND VDPWR VDPWR VGND _0626_ net56 net91 net104 dig_ctrl_inst.latch_mem_inst.RAM\[43\]\[6\]
+ sky130_fd_sc_hd__and4_1
X_2403_ VGND VDPWR VDPWR VGND clknet_leaf_6_clk _0011_ net146 dig_ctrl_inst.cpu_inst.port_o\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_153 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
X_1782_ VGND VDPWR VDPWR VGND _0491_ net62 net103 net131 dig_ctrl_inst.latch_mem_inst.RAM\[19\]\[3\]
+ sky130_fd_sc_hd__and4_1
X_2334_ VGND VDPWR VDPWR VGND _0086_ dig_ctrl_inst.spi_data_o\[7\] _0180_ dig_ctrl_inst.spi_data_o\[6\]
+ sky130_fd_sc_hd__mux2_1
X_2196_ VGND VDPWR VDPWR VGND _0884_ _0240_ _0885_ sky130_fd_sc_hd__xnor2_1
X_2265_ VGND VDPWR VDPWR VGND _0950_ _0236_ _0951_ sky130_fd_sc_hd__xnor2_1
X_1216_ VDPWR VGND VDPWR VGND _1064_ net254 net258 dig_ctrl_inst.cpu_inst.r3\[0\]
+ sky130_fd_sc_hd__and3_2
XFILLER_0_15_131 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_15_197 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xhold66 VGND VDPWR VDPWR VGND net348 dig_ctrl_inst.spi_data_i\[4\] sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 VGND VDPWR VDPWR VGND net326 dig_ctrl_inst.latch_mem_inst.wdata\[5\] sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 VGND VDPWR VDPWR VGND net370 dig_ctrl_inst.cpu_inst.r3\[3\] sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 VGND VDPWR VDPWR VGND net359 dig_ctrl_inst.cpu_inst.r1\[4\] sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 VGND VDPWR VDPWR VGND net381 dig_ctrl_inst.cpu_inst.r2\[3\] sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 VGND VDPWR VDPWR VGND net337 dig_ctrl_inst.spi_receiver_inst.synchronizer_spi_cs.pipe\[0\]
+ sky130_fd_sc_hd__dlygate4sd3_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[61\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[61\]\[4\] net210 dig_ctrl_inst.latch_mem_inst.gclk\[61\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[50\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[50\]\[2\] net228 dig_ctrl_inst.latch_mem_inst.gclk\[50\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_7_Left_85 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XANTENNA_8 VGND VDPWR VDPWR VGND _0674_ sky130_fd_sc_hd__diode_2
X_2050_ VDPWR VGND VDPWR VGND _1012_ dig_ctrl_inst.cpu_inst.instr\[5\] _0743_ net296
+ _1013_ sky130_fd_sc_hd__o211a_2
X_1834_ VGND VDPWR VDPWR VGND _1142_ dig_ctrl_inst.latch_mem_inst.RAM\[8\]\[4\] _0539_
+ _0540_ _0541_ _0542_ sky130_fd_sc_hd__a2111o_1
X_1903_ VDPWR VGND VDPWR VGND _0610_ net61 net109 dig_ctrl_inst.latch_mem_inst.RAM\[18\]\[5\]
+ sky130_fd_sc_hd__and3_2
X_1765_ VDPWR VGND VDPWR VGND _0474_ net67 net86 dig_ctrl_inst.latch_mem_inst.RAM\[24\]\[3\]
+ sky130_fd_sc_hd__and3_2
X_1696_ VGND VDPWR VDPWR VGND _0406_ net66 net91 net105 dig_ctrl_inst.latch_mem_inst.RAM\[27\]\[2\]
+ sky130_fd_sc_hd__and4_1
X_2317_ VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_receiver_inst.spi_sclk_delayed dig_ctrl_inst.spi_receiver_inst.spi_sclk_sync
+ dig_ctrl_inst.spi_receiver_inst.spi_cs_sync _0978_ sky130_fd_sc_hd__or3b_1
XFILLER_0_32_3 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_2248_ VGND VDPWR VDPWR VGND _0933_ _0935_ _0934_ sky130_fd_sc_hd__nand2_1
X_2179_ VGND VDPWR VDPWR VGND _0867_ _0869_ _0868_ sky130_fd_sc_hd__nand2_1
Xoutput23 VDPWR VGND VDPWR VGND port_ms_o[6] net23 sky130_fd_sc_hd__buf_2
Xoutput34 VDPWR VGND VDPWR VGND uo_out[6] net34 sky130_fd_sc_hd__buf_2
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[16\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[16\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[16\] clknet_leaf_15_clk sky130_fd_sc_hd__dlclkp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[54\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[54\]\[3\] net216 dig_ctrl_inst.latch_mem_inst.gclk\[54\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_5_109 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1481_ VGND VDPWR VDPWR VGND _0200_ dig_ctrl_inst.stb_dd _1039_ dig_ctrl_inst.stb_d
+ sky130_fd_sc_hd__mux2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[43\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[43\]\[1\] net234 dig_ctrl_inst.latch_mem_inst.gclk\[43\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_1_337 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1550_ VGND VDPWR VDPWR VGND net161 _0263_ net163 sky130_fd_sc_hd__and2b_1
X_2033_ VDPWR VGND VDPWR VGND _0720_ _0736_ _0735_ _0737_ _0738_ sky130_fd_sc_hd__or4_4
X_2102_ VDPWR VGND VDPWR VGND net164 _0747_ _0795_ dig_ctrl_inst.cpu_inst.data\[0\]
+ _0743_ sky130_fd_sc_hd__a22oi_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[34\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[34\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[34\] sky130_fd_sc_hd__clkbuf_4
X_1748_ VDPWR VGND VDPWR VGND _0136_ dig_ctrl_inst.latch_mem_inst.RAM\[18\]\[3\] _0121_
+ _0457_ dig_ctrl_inst.latch_mem_inst.RAM\[34\]\[3\] sky130_fd_sc_hd__a22o_1
X_1817_ VDPWR VGND VDPWR VGND _0525_ net84 net121 dig_ctrl_inst.latch_mem_inst.RAM\[10\]\[4\]
+ sky130_fd_sc_hd__and3_2
X_1679_ VGND VDPWR VDPWR VGND _0114_ dig_ctrl_inst.latch_mem_inst.RAM\[13\]\[1\] _0342_
+ _0343_ _0364_ _0390_ sky130_fd_sc_hd__a2111o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[20\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[20\]\[6\] net198 dig_ctrl_inst.latch_mem_inst.gclk\[20\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_64_29 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
Xdig_ctrl_inst.latch_mem_inst.gen_words\[58\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[58\]\[4\] net212 dig_ctrl_inst.latch_mem_inst.gclk\[58\]
+ sky130_fd_sc_hd__dlxtp_1
X_1602_ VGND VDPWR VDPWR VGND _0314_ net50 net112 dig_ctrl_inst.latch_mem_inst.RAM\[50\]\[0\]
+ _0129_ dig_ctrl_inst.latch_mem_inst.RAM\[26\]\[0\] sky130_fd_sc_hd__a32o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[47\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[47\]\[2\] net225 dig_ctrl_inst.latch_mem_inst.gclk\[47\]
+ sky130_fd_sc_hd__dlxtp_1
X_1464_ VGND VDPWR VDPWR VGND _0008_ _0192_ dig_ctrl_inst.spi_addr\[3\] _0193_ sky130_fd_sc_hd__mux2_1
X_1395_ VGND VDPWR VDPWR VGND _0153_ net102 net99 net42 sky130_fd_sc_hd__and3_4
X_1533_ VGND VDPWR VDPWR VGND net167 _0246_ net166 sky130_fd_sc_hd__nand2_1
Xfanout109 VDPWR VGND VDPWR VGND net109 net112 sky130_fd_sc_hd__buf_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[36\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[36\]\[0\] net246 dig_ctrl_inst.latch_mem_inst.gclk\[36\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_54_51 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_2016_ VDPWR VGND VDPWR VGND _0152_ dig_ctrl_inst.latch_mem_inst.RAM\[27\]\[7\] _0130_
+ _0721_ dig_ctrl_inst.latch_mem_inst.RAM\[54\]\[7\] sky130_fd_sc_hd__a22o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[2\].gen_latches\[6\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[2\]\[6\] net193 dig_ctrl_inst.latch_mem_inst.gclk\[2\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[24\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[24\]\[7\] net185 dig_ctrl_inst.latch_mem_inst.gclk\[24\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[13\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[13\]\[5\] net201 dig_ctrl_inst.latch_mem_inst.gclk\[13\]
+ sky130_fd_sc_hd__dlxtp_1
X_1180_ VGND VDPWR VDPWR VGND net297 net182 _1027_ _1028_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_20_Left_98 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_12_clk VGND VDPWR VDPWR VGND clknet_leaf_12_clk clknet_1_0__leaf_clk
+ sky130_fd_sc_hd__clkbuf_8
X_1516_ VGND VDPWR VDPWR VGND _0167_ net138 _0229_ sky130_fd_sc_hd__nor2_1
X_2496_ VGND VDPWR VDPWR VGND clknet_leaf_7_clk net343 net180 dig_ctrl_inst.stb_dd
+ sky130_fd_sc_hd__dfrtp_1
X_1447_ VDPWR VGND VDPWR VGND _0182_ _0181_ dig_ctrl_inst.spi_receiver_inst.spi_cnt\[1\]
+ dig_ctrl_inst.spi_receiver_inst.spi_cnt\[0\] sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[6\].gen_latches\[7\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[6\]\[7\] net187 dig_ctrl_inst.latch_mem_inst.gclk\[6\]
+ sky130_fd_sc_hd__dlxtp_1
X_1378_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[45\] net149 _0145_
+ sky130_fd_sc_hd__and2_1
Xfanout91 VGND VDPWR VDPWR VGND net92 net91 sky130_fd_sc_hd__clkbuf_2
Xfanout80 VDPWR VGND VDPWR VGND net80 net81 sky130_fd_sc_hd__buf_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[17\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[17\]\[6\] net195 dig_ctrl_inst.latch_mem_inst.gclk\[17\]
+ sky130_fd_sc_hd__dlxtp_1
X_2281_ VDPWR VGND VDPWR VGND _0966_ _0963_ _0949_ _0052_ sky130_fd_sc_hd__a21oi_1
X_1301_ VGND VDPWR VDPWR VGND net305 _1078_ _1048_ _1062_ _1093_ _1141_ sky130_fd_sc_hd__a2111oi_2
Xclkbuf_leaf_1_clk VGND VDPWR VDPWR VGND clknet_leaf_1_clk clknet_1_1__leaf_clk sky130_fd_sc_hd__clkbuf_8
X_2350_ VGND VDPWR VDPWR VGND _0100_ net33 _0987_ dig_ctrl_inst.cpu_inst.port_o\[5\]
+ sky130_fd_sc_hd__mux2_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[27\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[27\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[27\] sky130_fd_sc_hd__clkbuf_4
X_1232_ VDPWR VGND VDPWR VGND _1080_ dig_ctrl_inst.cpu_inst.r3\[1\] net255 net258
+ sky130_fd_sc_hd__and3_2
X_1163_ VGND VDPWR VDPWR VGND net258 _1011_ net254 sky130_fd_sc_hd__nand2b_2
X_1996_ VDPWR VGND VDPWR VGND _0148_ dig_ctrl_inst.latch_mem_inst.RAM\[47\]\[7\] _0146_
+ _0701_ dig_ctrl_inst.latch_mem_inst.RAM\[49\]\[7\] sky130_fd_sc_hd__a22o_1
XFILLER_0_51_96 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_62_3 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2479_ VGND VDPWR VDPWR VGND clknet_leaf_2_clk _0085_ net180 dig_ctrl_inst.spi_data_o\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload0 VGND VDPWR VDPWR VGND clkload0/Y clknet_1_0__leaf_clk sky130_fd_sc_hd__inv_8
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[23\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[23\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[23\] clknet_leaf_12_clk sky130_fd_sc_hd__dlclkp_1
X_1850_ VDPWR VGND VDPWR VGND _0556_ _0557_ _0555_ _0558_ sky130_fd_sc_hd__or3_1
XFILLER_0_21_44 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1781_ VGND VDPWR VDPWR VGND _0119_ dig_ctrl_inst.latch_mem_inst.RAM\[16\]\[3\] _0487_
+ _0488_ _0489_ _0490_ sky130_fd_sc_hd__a2111o_1
X_2333_ VGND VDPWR VDPWR VGND _0085_ dig_ctrl_inst.spi_data_o\[6\] _0180_ dig_ctrl_inst.spi_data_o\[5\]
+ sky130_fd_sc_hd__mux2_1
X_2402_ VGND VDPWR VDPWR VGND clknet_leaf_6_clk _0000_ net145 dig_ctrl_inst.cpu_inst.port_stb_o
+ sky130_fd_sc_hd__dfrtp_4
X_1215_ VGND VDPWR VDPWR VGND _1047_ net135 _1063_ sky130_fd_sc_hd__nor2_1
X_2195_ VGND VDPWR VDPWR VGND _0252_ _0864_ _0249_ _0884_ sky130_fd_sc_hd__o21a_1
X_2264_ VGND VDPWR VDPWR VGND _0228_ _0230_ _0927_ _0950_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_62_51 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_7_321 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_1979_ VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[0\]\[6\] _0671_ _0684_
+ _0288_ _0685_ sky130_fd_sc_hd__o22a_4
Xhold56 VGND VDPWR VDPWR VGND net338 dig_ctrl_inst.synchronizer_port_i_inst\[6\].pipe\[0\]
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 VGND VDPWR VDPWR VGND net327 dig_ctrl_inst.latch_mem_inst.wdata\[1\] sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 VGND VDPWR VDPWR VGND net349 dig_ctrl_inst.cpu_inst.prev_state\[1\] sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 VGND VDPWR VDPWR VGND net371 dig_ctrl_inst.cpu_inst.r2\[2\] sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 VGND VDPWR VDPWR VGND net360 dig_ctrl_inst.cpu_inst.r3\[0\] sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_51_Left_129 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XANTENNA_9 VGND VDPWR VDPWR VGND _1136_ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_60_Left_138 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[50\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[50\]\[6\] net192 dig_ctrl_inst.latch_mem_inst.gclk\[50\]
+ sky130_fd_sc_hd__dlxtp_1
X_1902_ VGND VDPWR VDPWR VGND _0609_ net42 net114 net131 dig_ctrl_inst.latch_mem_inst.RAM\[49\]\[5\]
+ sky130_fd_sc_hd__and4_1
X_1764_ VGND VDPWR VDPWR VGND _1145_ dig_ctrl_inst.latch_mem_inst.RAM\[11\]\[3\] _0470_
+ _0471_ _0472_ _0473_ sky130_fd_sc_hd__a2111o_1
X_1833_ VDPWR VGND VDPWR VGND _0541_ net65 net77 dig_ctrl_inst.latch_mem_inst.RAM\[28\]\[4\]
+ sky130_fd_sc_hd__and3_2
X_1695_ VGND VDPWR VDPWR VGND _0405_ net69 net107 net132 dig_ctrl_inst.latch_mem_inst.RAM\[19\]\[2\]
+ sky130_fd_sc_hd__and4_1
X_2316_ VGND VDPWR VDPWR VGND _0076_ _0975_ _0977_ net364 sky130_fd_sc_hd__mux2_1
X_2247_ VGND VDPWR VDPWR VGND net138 _0934_ _0911_ sky130_fd_sc_hd__nand2_1
X_2178_ VGND VDPWR VDPWR VGND net169 _0868_ _0842_ sky130_fd_sc_hd__nand2_1
Xoutput24 VDPWR VGND VDPWR VGND port_ms_o[7] net24 sky130_fd_sc_hd__buf_2
Xoutput35 VDPWR VGND VDPWR VGND uo_out[7] net35 sky130_fd_sc_hd__buf_2
XFILLER_0_11_190 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_19_Right_19 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[54\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[54\]\[7\] net189 dig_ctrl_inst.latch_mem_inst.gclk\[54\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_1_305 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_28_Right_28 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1480_ VDPWR VGND VDPWR VGND _0199_ _0198_ _0175_ _1023_ sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[43\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[43\]\[5\] net202 dig_ctrl_inst.latch_mem_inst.gclk\[43\]
+ sky130_fd_sc_hd__dlxtp_1
X_2032_ VGND VDPWR VDPWR VGND _0153_ dig_ctrl_inst.latch_mem_inst.RAM\[55\]\[7\] _0687_
+ _0695_ _0706_ _0737_ sky130_fd_sc_hd__a2111o_1
X_2101_ VGND VDPWR VDPWR VGND _0794_ _0791_ net158 _0786_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_37_Right_37 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[32\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[32\]\[3\] net217 dig_ctrl_inst.latch_mem_inst.gclk\[32\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_46_Right_46 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1747_ VGND VDPWR VDPWR VGND _0456_ net70 net73 dig_ctrl_inst.latch_mem_inst.RAM\[30\]\[3\]
+ _0156_ dig_ctrl_inst.latch_mem_inst.RAM\[59\]\[3\] sky130_fd_sc_hd__a32o_1
X_1816_ VGND VDPWR VDPWR VGND _0524_ net64 net104 net133 dig_ctrl_inst.latch_mem_inst.RAM\[19\]\[4\]
+ sky130_fd_sc_hd__and4_1
X_1678_ VGND VDPWR VDPWR VGND _0132_ dig_ctrl_inst.latch_mem_inst.RAM\[31\]\[1\] _0345_
+ _0346_ _0354_ _0389_ sky130_fd_sc_hd__a2111o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[21\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[21\]\[1\] net233 dig_ctrl_inst.latch_mem_inst.gclk\[21\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_55_Right_55 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_64_Right_64 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_73_Right_73 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[2\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[2\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[2\] clknet_leaf_12_clk sky130_fd_sc_hd__dlclkp_1
X_1601_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[31\]\[0\] _0132_ _0313_
+ _0277_ dig_ctrl_inst.latch_mem_inst.RAM\[4\]\[0\] _0312_ sky130_fd_sc_hd__a221o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[47\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[47\]\[6\] net197 dig_ctrl_inst.latch_mem_inst.gclk\[47\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[3\].gen_latches\[1\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[3\]\[1\] net238 dig_ctrl_inst.latch_mem_inst.gclk\[3\]
+ sky130_fd_sc_hd__dlxtp_1
X_1532_ VGND VDPWR VDPWR VGND _0237_ _0240_ _0244_ _0245_ sky130_fd_sc_hd__or3b_1
XFILLER_0_38_97 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1463_ VDPWR VGND VDPWR VGND _0193_ _0186_ _0191_ sky130_fd_sc_hd__and2_1
X_1394_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[54\] net42 net93
+ net148 sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[36\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[36\]\[4\] net208 dig_ctrl_inst.latch_mem_inst.gclk\[36\]
+ sky130_fd_sc_hd__dlxtp_1
X_2015_ VDPWR VGND VDPWR VGND _0705_ _0694_ _0693_ _0692_ _0720_ sky130_fd_sc_hd__or4_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[25\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[25\]\[2\] net224 dig_ctrl_inst.latch_mem_inst.gclk\[25\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_input_latches\[2\].n_latch VGND VDPWR VDPWR VGND
+ dig_ctrl_inst.latch_mem_inst.wdata\[2\] dig_ctrl_inst.data_out\[2\] clknet_leaf_8_clk
+ sky130_fd_sc_hd__dlxtn_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[14\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[14\]\[0\] net247 dig_ctrl_inst.latch_mem_inst.gclk\[14\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[28\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[28\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[28\] clknet_leaf_0_clk sky130_fd_sc_hd__dlclkp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[7\].gen_latches\[2\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[7\]\[2\] net229 dig_ctrl_inst.latch_mem_inst.gclk\[7\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_54_141 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_54_130 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_2495_ VGND VDPWR VDPWR VGND clknet_leaf_5_clk _0094_ net179 dig_ctrl_inst.spi_data_i\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[30\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[30\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[30\] clknet_leaf_0_clk sky130_fd_sc_hd__dlclkp_1
X_1515_ VDPWR VGND VDPWR VGND _0228_ _0167_ net138 sky130_fd_sc_hd__and2_1
X_1446_ VGND VDPWR VDPWR VGND _0180_ dig_ctrl_inst.spi_receiver_inst.spi_cnt\[0\]
+ _0002_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_65_51 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1377_ VDPWR VGND VDPWR VGND _0145_ net52 net80 net115 sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[29\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[29\]\[3\] net221 dig_ctrl_inst.latch_mem_inst.gclk\[29\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_5_271 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
Xdig_ctrl_inst.latch_mem_inst.gen_words\[18\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[18\]\[1\] net232 dig_ctrl_inst.latch_mem_inst.gclk\[18\]
+ sky130_fd_sc_hd__dlxtp_1
Xfanout92 VDPWR VGND VDPWR VGND _1140_ net92 sky130_fd_sc_hd__buf_4
Xfanout70 VDPWR VGND VDPWR VGND net70 net71 sky130_fd_sc_hd__buf_2
XFILLER_0_36_141 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
Xfanout81 VDPWR VGND VDPWR VGND net81 _1146_ sky130_fd_sc_hd__buf_2
X_2280_ VGND VDPWR VDPWR VGND _0965_ _0756_ _0964_ _0754_ _0966_ net41 sky130_fd_sc_hd__o221a_1
X_1231_ VGND VDPWR VDPWR VGND _1079_ _1026_ net182 _1027_ dig_ctrl_inst.cpu_inst.ip\[1\]
+ sky130_fd_sc_hd__o211a_1
X_1300_ VGND VDPWR VDPWR VGND net136 net135 _1140_ sky130_fd_sc_hd__nor2_1
X_1162_ VGND VDPWR VDPWR VGND net248 _1010_ dig_ctrl_inst.cpu_inst.cpu_state\[1\]
+ dig_ctrl_inst.cpu_inst.cpu_state\[2\] sky130_fd_sc_hd__nor3b_2
XFILLER_0_19_44 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_35_21 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_111 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_42_122 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
X_1995_ VDPWR VGND VDPWR VGND _0700_ net54 net96 dig_ctrl_inst.latch_mem_inst.RAM\[36\]\[7\]
+ sky130_fd_sc_hd__and3_2
X_2478_ VGND VDPWR VDPWR VGND clknet_leaf_4_clk _0084_ net172 dig_ctrl_inst.spi_data_o\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_3 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
X_1429_ VGND VDPWR VDPWR VGND net255 _0170_ dig_ctrl_inst.cpu_inst.r1\[7\] sky130_fd_sc_hd__and2b_1
Xclkload1 VGND VDPWR VDPWR VGND clkload1/Y clknet_leaf_10_clk sky130_fd_sc_hd__inv_16
Xfanout260 VDPWR VGND VDPWR VGND net261 net260 sky130_fd_sc_hd__buf_4
X_1780_ VDPWR VGND VDPWR VGND _0489_ net294 net121 dig_ctrl_inst.latch_mem_inst.RAM\[10\]\[3\]
+ sky130_fd_sc_hd__and3_2
X_2332_ VGND VDPWR VDPWR VGND _0084_ dig_ctrl_inst.spi_data_o\[5\] _0180_ dig_ctrl_inst.spi_data_o\[4\]
+ sky130_fd_sc_hd__mux2_1
X_2401_ VGND VDPWR VDPWR VGND clknet_leaf_4_clk _0010_ net176 dig_ctrl_inst.spi_addr\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_1214_ VGND VDPWR VDPWR VGND _1055_ _1061_ _1002_ _1062_ _1049_ dig_ctrl_inst.spi_addr\[2\]
+ sky130_fd_sc_hd__o32a_4
X_2194_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.r0\[4\] _0758_ _0883_ sky130_fd_sc_hd__nor2_1
X_2263_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.r0\[7\] net41 _0949_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_85 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_7_333 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[62\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[62\]\[3\] net221 dig_ctrl_inst.latch_mem_inst.gclk\[62\]
+ sky130_fd_sc_hd__dlxtp_1
X_1978_ VDPWR VGND VDPWR VGND _0683_ _0679_ _0674_ _0287_ _0684_ sky130_fd_sc_hd__or4_4
Xhold57 VGND VDPWR VDPWR VGND net339 dig_ctrl_inst.synchronizer_port_i_inst\[7\].pipe\[0\]
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 VGND VDPWR VDPWR VGND net328 dig_ctrl_inst.latch_mem_inst.wdata\[7\] sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 VGND VDPWR VDPWR VGND net350 dig_ctrl_inst.spi_data_i\[6\] sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 VGND VDPWR VDPWR VGND net361 dig_ctrl_inst.cpu_inst.r1\[6\] sky130_fd_sc_hd__dlygate4sd3_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[7\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[7\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[7\] clknet_leaf_1_clk sky130_fd_sc_hd__dlclkp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[51\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[51\]\[1\] net233 dig_ctrl_inst.latch_mem_inst.gclk\[51\]
+ sky130_fd_sc_hd__dlxtp_1
X_1901_ VGND VDPWR VDPWR VGND _0608_ net52 net90 net114 dig_ctrl_inst.latch_mem_inst.RAM\[41\]\[5\]
+ sky130_fd_sc_hd__and4_1
X_1832_ VDPWR VGND VDPWR VGND _0540_ net45 net96 dig_ctrl_inst.latch_mem_inst.RAM\[52\]\[4\]
+ sky130_fd_sc_hd__and3_2
X_1694_ VDPWR VGND VDPWR VGND _0404_ dig_ctrl_inst.latch_mem_inst.RAM\[43\]\[2\] _0143_
+ sky130_fd_sc_hd__and2_1
X_1763_ VGND VDPWR VDPWR VGND _0472_ net49 net106 net132 dig_ctrl_inst.latch_mem_inst.RAM\[51\]\[3\]
+ sky130_fd_sc_hd__and4_1
XFILLER_0_57_52 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2246_ VGND VDPWR VDPWR VGND _0933_ net138 _0911_ sky130_fd_sc_hd__or2_1
X_2315_ VGND VDPWR VDPWR VGND _0075_ _0974_ _0977_ net352 sky130_fd_sc_hd__mux2_1
X_2177_ VGND VDPWR VDPWR VGND _0867_ net169 _0842_ sky130_fd_sc_hd__or2_1
Xoutput25 VDPWR VGND VDPWR VGND uio_out[2] net25 sky130_fd_sc_hd__buf_2
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[59\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[59\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[59\] sky130_fd_sc_hd__clkbuf_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[55\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[55\]\[2\] net224 dig_ctrl_inst.latch_mem_inst.gclk\[55\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[44\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[44\]\[0\] net244 dig_ctrl_inst.latch_mem_inst.gclk\[44\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_1_317 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[35\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[35\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[35\] clknet_leaf_16_clk sky130_fd_sc_hd__dlclkp_1
X_2100_ VDPWR VGND VDPWR VGND _0793_ _1016_ _0745_ sky130_fd_sc_hd__or2_2
X_2031_ VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[11\]\[7\] _1145_ _0691_
+ _0698_ _0703_ _0736_ sky130_fd_sc_hd__a2111o_1
X_1815_ VGND VDPWR VDPWR VGND _0132_ dig_ctrl_inst.latch_mem_inst.RAM\[31\]\[4\] _0520_
+ _0521_ _0522_ _0523_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_32_209 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[32\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[32\]\[7\] net187 dig_ctrl_inst.latch_mem_inst.gclk\[32\]
+ sky130_fd_sc_hd__dlxtp_1
X_1746_ VDPWR VGND VDPWR VGND _0159_ dig_ctrl_inst.latch_mem_inst.RAM\[22\]\[3\] _0125_
+ _0455_ dig_ctrl_inst.latch_mem_inst.RAM\[62\]\[3\] sky130_fd_sc_hd__a22o_1
X_1677_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[15\]\[1\] _0117_ _0388_
+ _0143_ dig_ctrl_inst.latch_mem_inst.RAM\[43\]\[1\] _0367_ sky130_fd_sc_hd__a221o_1
X_2229_ VGND VDPWR VDPWR VGND _0917_ _0241_ _0243_ _0787_ _0914_ _0916_ sky130_fd_sc_hd__o311a_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[21\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[21\]\[5\] net202 dig_ctrl_inst.latch_mem_inst.gclk\[21\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[59\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[59\]\[3\] net222 dig_ctrl_inst.latch_mem_inst.gclk\[59\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[10\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[10\]\[3\] net217 dig_ctrl_inst.latch_mem_inst.gclk\[10\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_7_3 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[48\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[48\]\[1\] net236 dig_ctrl_inst.latch_mem_inst.gclk\[48\]
+ sky130_fd_sc_hd__dlxtp_1
X_1462_ VDPWR VGND VDPWR VGND _0007_ _0190_ _0192_ sky130_fd_sc_hd__and2_1
X_1600_ VGND VDPWR VDPWR VGND _0312_ net69 net74 dig_ctrl_inst.latch_mem_inst.RAM\[30\]\[0\]
+ _0142_ dig_ctrl_inst.latch_mem_inst.RAM\[42\]\[0\] sky130_fd_sc_hd__a32o_1
X_1531_ VGND VDPWR VDPWR VGND _0241_ _0243_ _0244_ sky130_fd_sc_hd__nor2_1
X_1393_ VDPWR VGND VDPWR VGND net94 net46 _0152_ sky130_fd_sc_hd__and2_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[3\].gen_latches\[5\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[3\]\[5\] net201 dig_ctrl_inst.latch_mem_inst.gclk\[3\]
+ sky130_fd_sc_hd__dlxtp_1
X_2014_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[8\]\[7\] _1142_ _0719_
+ _0142_ dig_ctrl_inst.latch_mem_inst.RAM\[42\]\[7\] _0718_ sky130_fd_sc_hd__a221o_1
XFILLER_0_49_139 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_49_117 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xhold110 VGND VDPWR VDPWR VGND net392 net18 sky130_fd_sc_hd__dlygate4sd3_1
X_1729_ VDPWR VGND VDPWR VGND _0436_ _0438_ _0437_ _0432_ _0439_ sky130_fd_sc_hd__or4_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[30\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[30\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[30\] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_13_297 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
Xdig_ctrl_inst.latch_mem_inst.gen_input_latches\[6\].n_latch VGND VDPWR VDPWR VGND
+ dig_ctrl_inst.latch_mem_inst.wdata\[6\] dig_ctrl_inst.data_out\[6\] clknet_leaf_8_clk
+ sky130_fd_sc_hd__dlxtn_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[25\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[25\]\[6\] net194 dig_ctrl_inst.latch_mem_inst.gclk\[25\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[14\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[14\]\[4\] net213 dig_ctrl_inst.latch_mem_inst.gclk\[14\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_51_337 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_24_23 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_54_153 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1445_ VDPWR VGND VDPWR VGND _0181_ _0180_ sky130_fd_sc_hd__inv_2
X_2494_ VGND VDPWR VDPWR VGND clknet_leaf_6_clk _0093_ net179 dig_ctrl_inst.spi_data_i\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[7\].gen_latches\[6\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[7\]\[6\] net198 dig_ctrl_inst.latch_mem_inst.gclk\[7\]
+ sky130_fd_sc_hd__dlxtp_1
X_1514_ VDPWR VGND VDPWR VGND _0227_ net265 net262 dig_ctrl_inst.cpu_inst.r0\[6\]
+ _0226_ _0225_ sky130_fd_sc_hd__o32a_1
XFILLER_0_65_63 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_1376_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[44\] net58 net78
+ net156 sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[29\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[29\]\[7\] net187 dig_ctrl_inst.latch_mem_inst.gclk\[29\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_28_109 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
Xdig_ctrl_inst.latch_mem_inst.gen_words\[18\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[18\]\[5\] net199 dig_ctrl_inst.latch_mem_inst.gclk\[18\]
+ sky130_fd_sc_hd__dlxtp_1
Xfanout82 VGND VDPWR VDPWR VGND _1146_ net82 sky130_fd_sc_hd__clkbuf_4
Xfanout60 VDPWR VGND VDPWR VGND _0133_ net60 sky130_fd_sc_hd__buf_6
Xfanout71 VGND VDPWR VDPWR VGND _0118_ net71 sky130_fd_sc_hd__clkbuf_2
Xfanout93 VDPWR VGND VDPWR VGND net93 net95 sky130_fd_sc_hd__buf_2
X_1161_ VGND VDPWR VDPWR VGND net248 dig_ctrl_inst.cpu_inst.cpu_state\[2\] _1009_
+ dig_ctrl_inst.cpu_inst.cpu_state\[1\] sky130_fd_sc_hd__nor3b_1
X_1230_ VDPWR VGND VDPWR VGND _1078_ dig_ctrl_inst.spi_addr\[0\] _1002_ sky130_fd_sc_hd__or2_2
X_1994_ VDPWR VGND VDPWR VGND _0699_ net55 net75 dig_ctrl_inst.latch_mem_inst.RAM\[46\]\[7\]
+ sky130_fd_sc_hd__and3_2
XFILLER_0_15_337 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2477_ VGND VDPWR VDPWR VGND clknet_leaf_4_clk _0083_ net172 dig_ctrl_inst.spi_data_o\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_1428_ VGND VDPWR VDPWR VGND net254 net258 _0169_ dig_ctrl_inst.cpu_inst.r2\[7\]
+ sky130_fd_sc_hd__and3b_1
X_1359_ VGND VDPWR VDPWR VGND _0137_ net131 net102 net51 sky130_fd_sc_hd__and3_4
Xclkload2 VGND VDPWR VDPWR VGND clkload2/Y clknet_leaf_11_clk sky130_fd_sc_hd__inv_12
Xfanout250 VGND VDPWR VDPWR VGND net251 net250 sky130_fd_sc_hd__clkbuf_2
Xfanout261 VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.arg1\[0\] net261 sky130_fd_sc_hd__clkbuf_2
X_2400_ VGND VDPWR VDPWR VGND clknet_leaf_4_clk _0009_ net176 dig_ctrl_inst.spi_addr\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_57 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
X_2262_ VDPWR VGND VDPWR VGND _0948_ _0943_ _0926_ _0051_ sky130_fd_sc_hd__a21oi_1
X_2331_ VGND VDPWR VDPWR VGND _0083_ dig_ctrl_inst.spi_data_o\[4\] _0180_ dig_ctrl_inst.spi_data_o\[3\]
+ sky130_fd_sc_hd__mux2_1
X_1213_ VDPWR VGND VDPWR VGND _1060_ _1039_ net249 _1061_ sky130_fd_sc_hd__a21o_1
X_2193_ VDPWR VGND VDPWR VGND _0882_ _0877_ _0858_ _0048_ sky130_fd_sc_hd__a21oi_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[42\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[42\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[42\] clknet_leaf_0_clk sky130_fd_sc_hd__dlclkp_1
X_1977_ VDPWR VGND VDPWR VGND _0682_ _0681_ _0680_ _0666_ _0683_ sky130_fd_sc_hd__or4_4
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[23\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[23\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[23\] sky130_fd_sc_hd__clkbuf_4
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[9\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[9\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[9\] sky130_fd_sc_hd__clkbuf_4
X_2529_ VGND VDPWR VDPWR VGND net25 dig_ctrl_inst.spi_miso_o sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_137 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xhold47 VGND VDPWR VDPWR VGND net329 dig_ctrl_inst.latch_mem_inst.wdata\[3\] sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 VGND VDPWR VDPWR VGND net351 dig_ctrl_inst.spi_data_i\[7\] sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 VGND VDPWR VDPWR VGND net340 dig_ctrl_inst.synchronizer_port_ms_i_inst.pipe\[0\]
+ sky130_fd_sc_hd__dlygate4sd3_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[62\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[62\]\[7\] net189 dig_ctrl_inst.latch_mem_inst.gclk\[62\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[51\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[51\]\[5\] net202 dig_ctrl_inst.latch_mem_inst.gclk\[51\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[40\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[40\]\[3\] net216 dig_ctrl_inst.latch_mem_inst.gclk\[40\]
+ sky130_fd_sc_hd__dlxtp_1
X_1831_ VDPWR VGND VDPWR VGND _0539_ net64 net72 dig_ctrl_inst.latch_mem_inst.RAM\[30\]\[4\]
+ sky130_fd_sc_hd__and3_2
X_1900_ VGND VDPWR VDPWR VGND _0135_ dig_ctrl_inst.latch_mem_inst.RAM\[33\]\[5\] _0604_
+ _0605_ _0606_ _0607_ sky130_fd_sc_hd__a2111o_1
X_1762_ VGND VDPWR VDPWR VGND _0471_ net59 net92 net119 dig_ctrl_inst.latch_mem_inst.RAM\[41\]\[3\]
+ sky130_fd_sc_hd__and4_1
X_1693_ VDPWR VGND VDPWR VGND _0403_ net78 net126 dig_ctrl_inst.latch_mem_inst.RAM\[12\]\[2\]
+ sky130_fd_sc_hd__and3_2
X_2314_ VGND VDPWR VDPWR VGND _0074_ _0973_ _0977_ net368 sky130_fd_sc_hd__mux2_1
X_2176_ VGND VDPWR VDPWR VGND _0864_ _0865_ _0866_ _0252_ sky130_fd_sc_hd__o21ai_1
X_2245_ VDPWR VGND VDPWR VGND net167 _0838_ _0932_ _0929_ _0931_ net170 sky130_fd_sc_hd__a221o_1
XFILLER_0_73_41 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xoutput26 VDPWR VGND VDPWR VGND uio_out[6] net26 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_1_Right_1 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[55\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[55\]\[6\] net197 dig_ctrl_inst.latch_mem_inst.gclk\[55\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[44\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[44\]\[4\] net209 dig_ctrl_inst.latch_mem_inst.gclk\[44\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_1_329 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
X_2030_ VGND VDPWR VDPWR VGND _0143_ dig_ctrl_inst.latch_mem_inst.RAM\[43\]\[7\] _0696_
+ _0697_ _0707_ _0735_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_43_77 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
Xdig_ctrl_inst.latch_mem_inst.gen_words\[33\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[33\]\[2\] net231 dig_ctrl_inst.latch_mem_inst.gclk\[33\]
+ sky130_fd_sc_hd__dlxtp_1
X_1745_ VDPWR VGND VDPWR VGND _0277_ dig_ctrl_inst.latch_mem_inst.RAM\[63\]\[3\] _0160_
+ _0454_ dig_ctrl_inst.latch_mem_inst.RAM\[4\]\[3\] sky130_fd_sc_hd__a22o_1
X_1814_ VDPWR VGND VDPWR VGND _0522_ net45 net76 dig_ctrl_inst.latch_mem_inst.RAM\[60\]\[4\]
+ sky130_fd_sc_hd__and3_2
XFILLER_0_68_85 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
Xdig_ctrl_inst.latch_mem_inst.gen_words\[22\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[22\]\[0\] net245 dig_ctrl_inst.latch_mem_inst.gclk\[22\]
+ sky130_fd_sc_hd__dlxtp_1
X_1676_ VGND VDPWR VDPWR VGND _0137_ dig_ctrl_inst.latch_mem_inst.RAM\[35\]\[1\] _0353_
+ _0356_ _0368_ _0387_ sky130_fd_sc_hd__a2111o_1
X_2228_ VDPWR VGND VDPWR VGND _0783_ net138 _0915_ _0916_ sky130_fd_sc_hd__a21oi_1
X_2159_ VDPWR VGND VDPWR VGND _0850_ _0247_ _0849_ _0248_ _0787_ sky130_fd_sc_hd__o2bb2a_1
XPHY_EDGE_ROW_39_Left_117 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[59\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[59\]\[7\] net188 dig_ctrl_inst.latch_mem_inst.gclk\[59\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[10\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[10\]\[7\] net185 dig_ctrl_inst.latch_mem_inst.gclk\[10\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_48_Left_126 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[4\].gen_latches\[0\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[4\]\[0\] net246 dig_ctrl_inst.latch_mem_inst.gclk\[4\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_57_Left_135 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[48\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[48\]\[5\] net201 dig_ctrl_inst.latch_mem_inst.gclk\[48\]
+ sky130_fd_sc_hd__dlxtp_1
X_1461_ VGND VDPWR VDPWR VGND _0192_ _1003_ _1096_ _0189_ _0184_ sky130_fd_sc_hd__o31a_1
X_1392_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[53\] net149 _0151_
+ sky130_fd_sc_hd__and2_1
X_1530_ VGND VDPWR VDPWR VGND _1103_ net160 _0243_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_66_Left_144 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2013_ VDPWR VGND VDPWR VGND _0156_ dig_ctrl_inst.latch_mem_inst.RAM\[19\]\[7\] _0122_
+ _0718_ dig_ctrl_inst.latch_mem_inst.RAM\[59\]\[7\] sky130_fd_sc_hd__a22o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[37\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[37\]\[3\] net217 dig_ctrl_inst.latch_mem_inst.gclk\[37\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[16\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[16\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[16\] sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_75_Left_153 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_15_clk VGND VDPWR VDPWR VGND clknet_leaf_15_clk clknet_1_0__leaf_clk
+ sky130_fd_sc_hd__clkbuf_8
Xhold100 VGND VDPWR VDPWR VGND net382 dig_ctrl_inst.spi_addr\[0\] sky130_fd_sc_hd__dlygate4sd3_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[26\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[26\]\[1\] net236 dig_ctrl_inst.latch_mem_inst.gclk\[26\]
+ sky130_fd_sc_hd__dlxtp_1
X_1728_ VGND VDPWR VDPWR VGND _0141_ dig_ctrl_inst.latch_mem_inst.RAM\[41\]\[2\] _0406_
+ _0408_ _0412_ _0438_ sky130_fd_sc_hd__a2111o_1
X_1659_ VDPWR VGND VDPWR VGND _0370_ net54 net76 dig_ctrl_inst.latch_mem_inst.RAM\[44\]\[1\]
+ sky130_fd_sc_hd__and3_2
XFILLER_0_0_181 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
X_2524__273 VGND VDPWR VDPWR VGND net273 _2524__273/HI sky130_fd_sc_hd__conb_1
XFILLER_0_39_151 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2531__277 VGND VDPWR VDPWR VGND net277 _2531__277/HI sky130_fd_sc_hd__conb_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[8\].gen_latches\[1\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[8\]\[1\] net235 dig_ctrl_inst.latch_mem_inst.gclk\[8\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_40_34 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[47\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[47\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[47\] clknet_leaf_18_clk sky130_fd_sc_hd__dlclkp_1
Xclkbuf_leaf_4_clk VGND VDPWR VDPWR VGND clknet_leaf_4_clk clknet_1_1__leaf_clk sky130_fd_sc_hd__clkbuf_8
X_2493_ VGND VDPWR VDPWR VGND clknet_leaf_6_clk _0092_ net179 dig_ctrl_inst.spi_data_i\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_1444_ VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_receiver_inst.spi_sclk_delayed _0180_
+ dig_ctrl_inst.spi_receiver_inst.spi_cs_sync dig_ctrl_inst.spi_receiver_inst.spi_sclk_sync
+ sky130_fd_sc_hd__or3b_4
X_1375_ VDPWR VGND VDPWR VGND _0144_ net78 net58 sky130_fd_sc_hd__and2_1
XFILLER_0_10_279 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_1513_ VDPWR VGND VDPWR VGND _0998_ dig_ctrl_inst.cpu_inst.r2\[6\] _0226_ dig_ctrl_inst.cpu_inst.r1\[6\]
+ _1022_ net299 sky130_fd_sc_hd__a221o_1
X_1159__1 VDPWR VGND VDPWR VGND net282 clknet_leaf_4_clk sky130_fd_sc_hd__inv_2
XFILLER_0_45_165 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_18_313 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[19\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[19\]\[0\] net244 dig_ctrl_inst.latch_mem_inst.gclk\[19\]
+ sky130_fd_sc_hd__dlxtp_1
Xfanout83 VDPWR VGND VDPWR VGND net83 net84 sky130_fd_sc_hd__buf_2
Xfanout50 VDPWR VGND VDPWR VGND _0147_ net50 sky130_fd_sc_hd__buf_4
Xfanout94 VGND VDPWR VDPWR VGND net94 net95 sky130_fd_sc_hd__buf_1
Xfanout72 VGND VDPWR VDPWR VGND net75 net72 sky130_fd_sc_hd__clkbuf_4
Xfanout61 VGND VDPWR VDPWR VGND net67 net61 sky130_fd_sc_hd__clkbuf_2
X_1160_ VGND VDPWR VDPWR VGND _1008_ _1002_ dig_ctrl_inst.spi_addr\[3\] sky130_fd_sc_hd__or2_1
X_1993_ VDPWR VGND VDPWR VGND _0698_ net48 net88 dig_ctrl_inst.latch_mem_inst.RAM\[56\]\[7\]
+ sky130_fd_sc_hd__and3_2
X_2476_ VGND VDPWR VDPWR VGND clknet_leaf_2_clk _0082_ net172 dig_ctrl_inst.spi_data_o\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_1427_ VDPWR VGND VDPWR VGND _0168_ dig_ctrl_inst.cpu_inst.r3\[7\] net255 net258
+ sky130_fd_sc_hd__and3_2
X_1358_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[34\] net51 net109
+ net148 sky130_fd_sc_hd__and3_2
X_1289_ VGND VDPWR VDPWR VGND _1134_ net304 _1078_ _1093_ sky130_fd_sc_hd__and3_4
Xclkload3 VGND VDPWR VDPWR VGND clknet_leaf_12_clk clkload3/Y sky130_fd_sc_hd__clkinv_8
Xfanout240 VGND VDPWR VDPWR VGND net241 net240 sky130_fd_sc_hd__clkbuf_2
Xfanout251 VGND VDPWR VDPWR VGND dig_ctrl_inst.mode_sync net251 sky130_fd_sc_hd__clkbuf_2
Xfanout262 VDPWR VGND VDPWR VGND net264 net262 sky130_fd_sc_hd__buf_4
X_2330_ VGND VDPWR VDPWR VGND _0082_ dig_ctrl_inst.spi_data_o\[3\] _0180_ dig_ctrl_inst.spi_data_o\[2\]
+ sky130_fd_sc_hd__mux2_1
X_1212_ VGND VDPWR VDPWR VGND net300 _1056_ _1057_ _1058_ _1059_ _1060_ sky130_fd_sc_hd__o41a_2
X_2192_ VGND VDPWR VDPWR VGND _0881_ _0756_ _0880_ _0754_ _0882_ net41 sky130_fd_sc_hd__o221a_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[62\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[62\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[62\] sky130_fd_sc_hd__clkbuf_4
X_2261_ VGND VDPWR VDPWR VGND _0947_ _0756_ _0946_ _0754_ _0948_ net41 sky130_fd_sc_hd__o221a_1
XFILLER_0_47_205 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[63\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[63\]\[2\] net226 dig_ctrl_inst.latch_mem_inst.gclk\[63\]
+ sky130_fd_sc_hd__dlxtp_1
X_1976_ VGND VDPWR VDPWR VGND _0141_ dig_ctrl_inst.latch_mem_inst.RAM\[41\]\[6\] _0626_
+ _0627_ _0629_ _0682_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_15_146 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2528_ VDPWR VGND VDPWR VGND uio_out[1] net275 sky130_fd_sc_hd__buf_2
Xhold48 VGND VDPWR VDPWR VGND net330 dig_ctrl_inst.synchronizer_port_i_inst\[3\].pipe\[0\]
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 VGND VDPWR VDPWR VGND net341 dig_ctrl_inst.synchronizer_port_i_inst\[0\].pipe\[0\]
+ sky130_fd_sc_hd__dlygate4sd3_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[52\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[52\]\[0\] net241 dig_ctrl_inst.latch_mem_inst.gclk\[52\]
+ sky130_fd_sc_hd__dlxtp_1
X_2459_ VGND VDPWR VDPWR VGND clknet_leaf_11_clk _0067_ net142 dig_ctrl_inst.cpu_inst.r2\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[40\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[40\]\[7\] net185 dig_ctrl_inst.latch_mem_inst.gclk\[40\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_16_69 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1761_ VGND VDPWR VDPWR VGND _0470_ net101 net106 net126 dig_ctrl_inst.latch_mem_inst.RAM\[7\]\[3\]
+ sky130_fd_sc_hd__and4_1
X_1830_ VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[57\]\[4\] _0154_ _0535_
+ _0536_ _0537_ _0538_ sky130_fd_sc_hd__a2111o_1
X_1692_ VDPWR VGND VDPWR VGND _0402_ net50 net88 dig_ctrl_inst.latch_mem_inst.RAM\[56\]\[2\]
+ sky130_fd_sc_hd__and3_2
X_2313_ VGND VDPWR VDPWR VGND _0073_ _0972_ _0977_ net376 sky130_fd_sc_hd__mux2_1
X_2175_ VDPWR VGND VDPWR VGND _0864_ _0252_ _0788_ _0865_ sky130_fd_sc_hd__a21oi_1
X_2244_ VDPWR VGND VDPWR VGND _0931_ _0930_ _0886_ _0840_ sky130_fd_sc_hd__and3_2
XPHY_EDGE_ROW_11_Left_89 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[56\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[56\]\[1\] net238 dig_ctrl_inst.latch_mem_inst.gclk\[56\]
+ sky130_fd_sc_hd__dlxtp_1
X_1959_ VGND VDPWR VDPWR VGND _0138_ dig_ctrl_inst.latch_mem_inst.RAM\[37\]\[6\] _0624_
+ _0647_ _0659_ _0665_ sky130_fd_sc_hd__a2111o_1
Xoutput27 VDPWR VGND VDPWR VGND uio_out[7] net27 sky130_fd_sc_hd__buf_2
Xoutput16 VGND VDPWR VDPWR VGND clk_o net16 sky130_fd_sc_hd__clkbuf_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[0\].gen_latches\[3\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[0\]\[3\] net218 dig_ctrl_inst.latch_mem_inst.gclk\[0\]
+ sky130_fd_sc_hd__dlxtp_1
Xclkbuf_0_clk VGND VDPWR VDPWR VGND clk clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_43_89 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
Xdig_ctrl_inst.latch_mem_inst.gen_words\[33\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[33\]\[6\] net192 dig_ctrl_inst.latch_mem_inst.gclk\[33\]
+ sky130_fd_sc_hd__dlxtp_1
X_1744_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[14\]\[3\] _0116_ _0453_
+ _0279_ dig_ctrl_inst.latch_mem_inst.RAM\[6\]\[3\] _0452_ sky130_fd_sc_hd__a221o_1
X_1813_ VDPWR VGND VDPWR VGND _0521_ net54 net76 dig_ctrl_inst.latch_mem_inst.RAM\[44\]\[4\]
+ sky130_fd_sc_hd__and3_2
XFILLER_0_4_179 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[22\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[22\]\[4\] net212 dig_ctrl_inst.latch_mem_inst.gclk\[22\]
+ sky130_fd_sc_hd__dlxtp_1
X_1675_ VDPWR VGND VDPWR VGND _0380_ _0385_ _0381_ _0379_ _0386_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_15_Right_15 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[54\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[54\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[54\] clknet_leaf_16_clk sky130_fd_sc_hd__dlclkp_1
XFILLER_0_23_3 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
X_2158_ VGND VDPWR VDPWR VGND _0849_ _0790_ net167 _0785_ sky130_fd_sc_hd__a21bo_1
X_2089_ VGND VDPWR VDPWR VGND _0782_ net171 _0781_ net168 _0774_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_24_Right_24 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2227_ VDPWR VGND VDPWR VGND _0825_ dig_ctrl_inst.cpu_inst.data\[5\] _0743_ _0915_
+ net159 sky130_fd_sc_hd__a22o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[11\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[11\]\[2\] net229 dig_ctrl_inst.latch_mem_inst.gclk\[11\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_33_Right_33 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[49\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[49\]\[0\] net244 dig_ctrl_inst.latch_mem_inst.gclk\[49\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_42_Right_42 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_51_Right_51 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[4\].gen_latches\[4\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[4\]\[4\] net213 dig_ctrl_inst.latch_mem_inst.gclk\[4\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[55\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[55\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[55\] sky130_fd_sc_hd__clkbuf_4
X_1460_ VGND VDPWR VDPWR VGND _1003_ _0189_ _0191_ sky130_fd_sc_hd__nor2_1
X_1391_ VDPWR VGND VDPWR VGND _0151_ net45 net100 net117 sky130_fd_sc_hd__and3_2
X_2012_ VDPWR VGND VDPWR VGND _0715_ _0716_ _0714_ _0717_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_60_Right_60 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[37\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[37\]\[7\] net186 dig_ctrl_inst.latch_mem_inst.gclk\[37\]
+ sky130_fd_sc_hd__dlxtp_1
X_1727_ VGND VDPWR VDPWR VGND _0139_ dig_ctrl_inst.latch_mem_inst.RAM\[39\]\[2\] _0403_
+ _0407_ _0409_ _0437_ sky130_fd_sc_hd__a2111o_1
Xhold101 VGND VDPWR VDPWR VGND net383 net23 sky130_fd_sc_hd__dlygate4sd3_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[26\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[26\]\[5\] net203 dig_ctrl_inst.latch_mem_inst.gclk\[26\]
+ sky130_fd_sc_hd__dlxtp_1
X_1658_ VDPWR VGND VDPWR VGND _0369_ net55 net128 dig_ctrl_inst.latch_mem_inst.RAM\[32\]\[1\]
+ sky130_fd_sc_hd__and3_2
X_1589_ VDPWR VGND VDPWR VGND _0301_ net74 net123 dig_ctrl_inst.latch_mem_inst.RAM\[14\]\[0\]
+ sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[15\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[15\]\[3\] net222 dig_ctrl_inst.latch_mem_inst.gclk\[15\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_14_Left_92 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[8\].gen_latches\[5\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[8\]\[5\] net204 dig_ctrl_inst.latch_mem_inst.gclk\[8\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_40_24 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2492_ VGND VDPWR VDPWR VGND clknet_leaf_4_clk _0091_ net179 dig_ctrl_inst.spi_data_i\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_57 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1512_ VDPWR VGND VDPWR VGND _0225_ dig_ctrl_inst.cpu_inst.r3\[6\] net262 net265
+ sky130_fd_sc_hd__and3_2
X_1443_ VDPWR VGND VDPWR VGND dig_ctrl_inst.cpu_inst.stb_o _0177_ _0178_ _0179_ _1027_
+ _1039_ sky130_fd_sc_hd__o32a_1
X_1374_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[43\] net152 _0143_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_65_87 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_45_144 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[19\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[19\]\[4\] net208 dig_ctrl_inst.latch_mem_inst.gclk\[19\]
+ sky130_fd_sc_hd__dlxtp_1
Xfanout73 VDPWR VGND VDPWR VGND net73 net74 sky130_fd_sc_hd__buf_2
Xfanout51 VDPWR VGND VDPWR VGND net53 net51 sky130_fd_sc_hd__buf_4
Xfanout62 VGND VDPWR VDPWR VGND net63 net62 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_51_125 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
Xfanout84 VDPWR VGND VDPWR VGND _1144_ net84 sky130_fd_sc_hd__buf_4
Xfanout95 VDPWR VGND VDPWR VGND _1138_ net95 sky130_fd_sc_hd__buf_4
XFILLER_0_24_339 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_35_57 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xclkload10 VDPWR VGND VDPWR VGND clknet_leaf_3_clk clkload10/Y sky130_fd_sc_hd__clkinv_4
X_1992_ VDPWR VGND VDPWR VGND _0697_ net64 net111 dig_ctrl_inst.latch_mem_inst.RAM\[18\]\[7\]
+ sky130_fd_sc_hd__and3_2
X_2475_ VGND VDPWR VDPWR VGND clknet_leaf_4_clk _0081_ net172 dig_ctrl_inst.spi_data_o\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_1426_ VDPWR VGND VDPWR VGND _0162_ net250 dig_ctrl_inst.spi_data_o\[6\] dig_ctrl_inst.data_out\[6\]
+ _0167_ sky130_fd_sc_hd__a22o_1
X_1357_ VDPWR VGND VDPWR VGND _0136_ net111 net58 sky130_fd_sc_hd__and2_1
X_1288_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[2\] net109 net120
+ net150 sky130_fd_sc_hd__and3_2
XFILLER_0_58_291 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xclkload4 VDPWR VGND VDPWR VGND clknet_leaf_13_clk clkload4/Y sky130_fd_sc_hd__clkinv_4
Xfanout263 VDPWR VGND VDPWR VGND net264 net263 sky130_fd_sc_hd__buf_6
Xfanout230 VGND VDPWR VDPWR VGND net231 net230 sky130_fd_sc_hd__clkbuf_2
Xfanout241 VGND VDPWR VDPWR VGND net242 net241 sky130_fd_sc_hd__clkbuf_2
Xfanout252 VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.instr\[5\] net252 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_21_15 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[48\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[48\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[48\] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_12_309 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
X_2191_ VDPWR VGND VDPWR VGND dig_ctrl_inst.spi_data_o\[3\] _0804_ _0881_ dig_ctrl_inst.synchronizer_port_i_inst\[3\].out
+ _0802_ sky130_fd_sc_hd__a22oi_1
X_1211_ VDPWR VGND VDPWR VGND net263 dig_ctrl_inst.cpu_inst.r0\[2\] net268 _1059_
+ sky130_fd_sc_hd__or3_1
X_2260_ VDPWR VGND VDPWR VGND dig_ctrl_inst.spi_data_o\[6\] _0804_ _0947_ dig_ctrl_inst.synchronizer_port_i_inst\[6\].out
+ _0802_ sky130_fd_sc_hd__a22oi_2
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[59\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[59\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[59\] clknet_leaf_0_clk sky130_fd_sc_hd__dlclkp_1
XFILLER_0_62_66 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
Xdig_ctrl_inst.latch_mem_inst.gen_words\[63\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[63\]\[6\] net194 dig_ctrl_inst.latch_mem_inst.gclk\[63\]
+ sky130_fd_sc_hd__dlxtp_1
X_1975_ VGND VDPWR VDPWR VGND _0149_ dig_ctrl_inst.latch_mem_inst.RAM\[51\]\[6\] _0628_
+ _0631_ _0653_ _0681_ sky130_fd_sc_hd__a2111o_1
X_2458_ VGND VDPWR VDPWR VGND clknet_leaf_7_clk _0066_ net143 dig_ctrl_inst.cpu_inst.r2\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_2527_ VDPWR VGND VDPWR VGND uio_out[0] net274 sky130_fd_sc_hd__buf_2
X_1409_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[62\] net48 net73
+ net153 sky130_fd_sc_hd__and3_2
X_2389_ VGND VDPWR VDPWR VGND clknet_leaf_4_clk net334 net172 dig_ctrl_inst.synchronizer_port_i_inst\[2\].out
+ sky130_fd_sc_hd__dfrtp_1
Xhold49 VGND VDPWR VDPWR VGND net331 dig_ctrl_inst.synchronizer_port_i_inst\[5\].pipe\[0\]
+ sky130_fd_sc_hd__dlygate4sd3_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[52\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[52\]\[4\] net209 dig_ctrl_inst.latch_mem_inst.gclk\[52\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[61\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[61\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[61\] clknet_leaf_15_clk sky130_fd_sc_hd__dlclkp_1
XFILLER_0_21_106 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
Xdig_ctrl_inst.latch_mem_inst.gen_words\[41\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[41\]\[2\] net225 dig_ctrl_inst.latch_mem_inst.gclk\[41\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[30\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[30\]\[0\] net244 dig_ctrl_inst.latch_mem_inst.gclk\[30\]
+ sky130_fd_sc_hd__dlxtp_1
X_1691_ VGND VDPWR VDPWR VGND _0401_ net82 net106 net127 dig_ctrl_inst.latch_mem_inst.RAM\[15\]\[2\]
+ sky130_fd_sc_hd__and4_1
XFILLER_0_52_253 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1760_ VDPWR VGND VDPWR VGND _0467_ _0468_ _0466_ _0469_ sky130_fd_sc_hd__or3_1
XFILLER_0_4_328 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_2_Left_80 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2312_ VGND VDPWR VDPWR VGND _0072_ _0971_ _0977_ net370 sky130_fd_sc_hd__mux2_1
X_2243_ VGND VDPWR VDPWR VGND _0930_ _0770_ _0775_ net158 _0778_ sky130_fd_sc_hd__a211o_1
X_2174_ VGND VDPWR VDPWR VGND _0248_ _0852_ _0246_ _0864_ sky130_fd_sc_hd__o21a_1
X_1889_ VDPWR VGND VDPWR VGND _0149_ dig_ctrl_inst.latch_mem_inst.RAM\[43\]\[5\] _0143_
+ _0596_ dig_ctrl_inst.latch_mem_inst.RAM\[51\]\[5\] sky130_fd_sc_hd__a22o_1
Xoutput28 VDPWR VGND VDPWR VGND uo_out[0] net28 sky130_fd_sc_hd__buf_2
Xoutput17 VDPWR VGND VDPWR VGND port_ms_o[0] net17 sky130_fd_sc_hd__buf_2
X_1958_ VDPWR VGND VDPWR VGND _0652_ _0655_ _0654_ _0640_ _0664_ sky130_fd_sc_hd__or4_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[56\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[56\]\[5\] net204 dig_ctrl_inst.latch_mem_inst.gclk\[56\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[5\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[5\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[5\] sky130_fd_sc_hd__clkbuf_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[45\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[45\]\[3\] net219 dig_ctrl_inst.latch_mem_inst.gclk\[45\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[34\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[34\]\[1\] net233 dig_ctrl_inst.latch_mem_inst.gclk\[34\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[0\].gen_latches\[7\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[0\]\[7\] net190 dig_ctrl_inst.latch_mem_inst.gclk\[0\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_27_69 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1743_ VDPWR VGND VDPWR VGND _0123_ dig_ctrl_inst.latch_mem_inst.RAM\[1\]\[3\] _1130_
+ _0452_ dig_ctrl_inst.latch_mem_inst.RAM\[20\]\[3\] sky130_fd_sc_hd__a22o_1
X_1812_ VDPWR VGND VDPWR VGND _0520_ net64 net129 dig_ctrl_inst.latch_mem_inst.RAM\[16\]\[4\]
+ sky130_fd_sc_hd__and3_2
X_1674_ VGND VDPWR VDPWR VGND _0154_ dig_ctrl_inst.latch_mem_inst.RAM\[57\]\[1\] _0355_
+ _0363_ _0366_ _0385_ sky130_fd_sc_hd__a2111o_1
X_2226_ VGND VDPWR VDPWR VGND _0793_ _0242_ _0785_ _0243_ _0914_ _0913_ sky130_fd_sc_hd__o221a_1
X_2157_ VGND VDPWR VDPWR VGND _0847_ _0246_ _0793_ _0848_ sky130_fd_sc_hd__o21ba_1
X_2088_ VGND VDPWR VDPWR VGND _0765_ _0777_ _0768_ _0780_ _0781_ sky130_fd_sc_hd__o22a_1
XFILLER_0_16_253 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_16_231 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[11\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[11\]\[6\] net195 dig_ctrl_inst.latch_mem_inst.gclk\[11\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[49\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[49\]\[4\] net212 dig_ctrl_inst.latch_mem_inst.gclk\[49\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[38\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[38\]\[2\] net228 dig_ctrl_inst.latch_mem_inst.gclk\[38\]
+ sky130_fd_sc_hd__dlxtp_1
X_1390_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[52\] net43 net96
+ net151 sky130_fd_sc_hd__and3_2
X_2011_ VDPWR VGND VDPWR VGND _0117_ dig_ctrl_inst.latch_mem_inst.RAM\[7\]\[7\] _1139_
+ _0716_ dig_ctrl_inst.latch_mem_inst.RAM\[15\]\[7\] sky130_fd_sc_hd__a22o_1
XFILLER_0_49_109 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[27\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[27\]\[0\] net241 dig_ctrl_inst.latch_mem_inst.gclk\[27\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_70_99 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_70_11 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1726_ VGND VDPWR VDPWR VGND _1145_ dig_ctrl_inst.latch_mem_inst.RAM\[11\]\[2\] _0399_
+ _0401_ _0410_ _0436_ sky130_fd_sc_hd__a2111o_1
X_1657_ VDPWR VGND VDPWR VGND _0368_ net86 net121 dig_ctrl_inst.latch_mem_inst.RAM\[8\]\[1\]
+ sky130_fd_sc_hd__and3_2
XFILLER_0_13_289 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1588_ VDPWR VGND VDPWR VGND _0300_ net45 net130 dig_ctrl_inst.latch_mem_inst.RAM\[48\]\[0\]
+ sky130_fd_sc_hd__and3_2
Xhold102 VGND VDPWR VDPWR VGND net384 dig_ctrl_inst.cpu_inst.r2\[7\] sky130_fd_sc_hd__dlygate4sd3_1
X_2209_ VGND VDPWR VDPWR VGND _0898_ _0239_ _0785_ _0895_ _0897_ sky130_fd_sc_hd__o211a_1
XFILLER_0_48_175 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
Xdig_ctrl_inst.latch_mem_inst.gen_words\[15\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[15\]\[7\] net189 dig_ctrl_inst.latch_mem_inst.gclk\[15\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[9\].gen_latches\[0\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[9\]\[0\] net241 dig_ctrl_inst.latch_mem_inst.gclk\[9\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_5_3 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_27_337 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2491_ VGND VDPWR VDPWR VGND clknet_leaf_5_clk _0090_ net178 dig_ctrl_inst.spi_data_i\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_1442_ VDPWR VGND VDPWR VGND dig_ctrl_inst.cpu_inst.cpu_state\[1\] _0179_ dig_ctrl_inst.cpu_inst.prev_state\[1\]
+ sky130_fd_sc_hd__xor2_1
X_1511_ VDPWR VGND VDPWR VGND _0024_ _1006_ _0220_ _0204_ _0224_ sky130_fd_sc_hd__o2bb2a_1
X_1373_ VDPWR VGND VDPWR VGND _0143_ net59 net92 net108 sky130_fd_sc_hd__and3_2
XFILLER_0_14_81 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[12\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[12\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[12\] sky130_fd_sc_hd__clkbuf_4
X_1709_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[1\]\[2\] _1130_ _0419_
+ _0160_ dig_ctrl_inst.latch_mem_inst.RAM\[63\]\[2\] _0418_ sky130_fd_sc_hd__a221o_1
Xfanout41 VDPWR VGND VDPWR VGND net41 _0758_ sky130_fd_sc_hd__buf_2
Xfanout74 VDPWR VGND VDPWR VGND net75 net74 sky130_fd_sc_hd__buf_4
Xfanout96 VDPWR VGND VDPWR VGND net96 net98 sky130_fd_sc_hd__buf_2
Xfanout63 VGND VDPWR VDPWR VGND net67 net63 sky130_fd_sc_hd__clkbuf_2
Xfanout52 VGND VDPWR VDPWR VGND net53 net52 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_51_137 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
Xdig_ctrl_inst.latch_mem_inst.gen_words\[60\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[60\]\[0\] net244 dig_ctrl_inst.latch_mem_inst.gclk\[60\]
+ sky130_fd_sc_hd__dlxtp_1
Xclkload11 VGND VDPWR VDPWR VGND clknet_leaf_4_clk clkload11/Y sky130_fd_sc_hd__bufinv_16
X_1991_ VDPWR VGND VDPWR VGND _0696_ net64 net130 dig_ctrl_inst.latch_mem_inst.RAM\[16\]\[7\]
+ sky130_fd_sc_hd__and3_2
X_2474_ VGND VDPWR VDPWR VGND clknet_leaf_4_clk _0080_ net172 dig_ctrl_inst.spi_data_o\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_1425_ VGND VDPWR VDPWR VGND _0167_ _0166_ _0165_ _0164_ _0163_ _1018_ sky130_fd_sc_hd__o41a_4
X_1356_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[33\] net150 _0135_
+ sky130_fd_sc_hd__and2_1
X_1287_ VDPWR VGND VDPWR VGND net120 net110 _1133_ sky130_fd_sc_hd__and2_2
Xclkload5 VGND VDPWR VDPWR VGND clkload5/Y clknet_leaf_15_clk sky130_fd_sc_hd__inv_8
Xfanout231 VDPWR VGND VDPWR VGND net231 net324 sky130_fd_sc_hd__buf_2
Xfanout264 VDPWR VGND VDPWR VGND dig_ctrl_inst.cpu_inst.arg0\[1\] net264 sky130_fd_sc_hd__buf_4
Xfanout220 VGND VDPWR VDPWR VGND net221 net220 sky130_fd_sc_hd__clkbuf_2
Xfanout242 VDPWR VGND VDPWR VGND net242 net247 sky130_fd_sc_hd__buf_2
Xfanout253 VDPWR VGND VDPWR VGND dig_ctrl_inst.cpu_inst.instr\[4\] net253 sky130_fd_sc_hd__buf_4
XFILLER_0_21_27 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_2190_ VGND VDPWR VDPWR VGND _0878_ _0879_ _0880_ sky130_fd_sc_hd__nand2b_1
X_1210_ VGND VDPWR VDPWR VGND net263 _1058_ dig_ctrl_inst.cpu_inst.r1\[2\] sky130_fd_sc_hd__and2b_1
XFILLER_0_62_12 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_1_15 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_78 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
X_1974_ VGND VDPWR VDPWR VGND _0151_ dig_ctrl_inst.latch_mem_inst.RAM\[53\]\[6\] _0634_
+ _0645_ _0651_ _0680_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_7_337 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2388_ VGND VDPWR VDPWR VGND clknet_leaf_4_clk net5 net174 dig_ctrl_inst.synchronizer_port_i_inst\[2\].pipe\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_2457_ VGND VDPWR VDPWR VGND clknet_leaf_7_clk _0065_ net143 dig_ctrl_inst.cpu_inst.r2\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_1408_ VDPWR VGND VDPWR VGND net73 net49 _0159_ sky130_fd_sc_hd__and2_2
X_2526_ VDPWR VGND VDPWR VGND uio_oe[7] net281 sky130_fd_sc_hd__buf_2
XFILLER_0_46_3 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_1339_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[24\] net67 net86
+ net149 sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[41\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[41\]\[6\] net193 dig_ctrl_inst.latch_mem_inst.gclk\[41\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[30\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[30\]\[4\] net209 dig_ctrl_inst.latch_mem_inst.gclk\[30\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_32_15 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1690_ VDPWR VGND VDPWR VGND _0400_ net58 net95 dig_ctrl_inst.latch_mem_inst.RAM\[38\]\[2\]
+ sky130_fd_sc_hd__and3_2
X_2311_ VGND VDPWR VDPWR VGND _0071_ _0970_ _0977_ net373 sky130_fd_sc_hd__mux2_1
X_2242_ VGND VDPWR VDPWR VGND _0929_ _0836_ _0887_ sky130_fd_sc_hd__or2_1
X_2173_ VGND VDPWR VDPWR VGND net170 _0862_ _0772_ _0860_ _0861_ _0863_ sky130_fd_sc_hd__a311o_1
X_1957_ VDPWR VGND VDPWR VGND _0157_ dig_ctrl_inst.latch_mem_inst.RAM\[7\]\[6\] _1139_
+ _0663_ dig_ctrl_inst.latch_mem_inst.RAM\[60\]\[6\] sky130_fd_sc_hd__a22o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[57\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[57\]\[0\] net245 dig_ctrl_inst.latch_mem_inst.gclk\[57\]
+ sky130_fd_sc_hd__dlxtp_1
X_2509_ VGND VDPWR VDPWR VGND clknet_leaf_5_clk _0106_ net178 net20 sky130_fd_sc_hd__dfrtp_1
Xoutput18 VDPWR VGND VDPWR VGND port_ms_o[1] net18 sky130_fd_sc_hd__buf_2
Xoutput29 VDPWR VGND VDPWR VGND uo_out[1] net29 sky130_fd_sc_hd__buf_2
X_1888_ VDPWR VGND VDPWR VGND _0124_ dig_ctrl_inst.latch_mem_inst.RAM\[17\]\[5\] _0120_
+ _0595_ dig_ctrl_inst.latch_mem_inst.RAM\[21\]\[5\] sky130_fd_sc_hd__a22o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[1\].gen_latches\[2\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[1\]\[2\] net226 dig_ctrl_inst.latch_mem_inst.gclk\[1\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[45\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[45\]\[7\] net184 dig_ctrl_inst.latch_mem_inst.gclk\[45\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[34\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[34\]\[5\] net199 dig_ctrl_inst.latch_mem_inst.gclk\[34\]
+ sky130_fd_sc_hd__dlxtp_1
X_1811_ VDPWR VGND VDPWR VGND _0508_ _0518_ _0511_ _0287_ _0519_ sky130_fd_sc_hd__or4_1
XFILLER_0_25_210 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1742_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[3\]\[3\] _1135_ _0451_
+ _0154_ dig_ctrl_inst.latch_mem_inst.RAM\[57\]\[3\] _0450_ sky130_fd_sc_hd__a221o_1
X_1673_ VDPWR VGND VDPWR VGND _0376_ _0383_ _0382_ _0374_ _0384_ sky130_fd_sc_hd__or4_1
XFILLER_0_0_321 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
Xdig_ctrl_inst.latch_mem_inst.gen_words\[23\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[23\]\[3\] net215 dig_ctrl_inst.latch_mem_inst.gclk\[23\]
+ sky130_fd_sc_hd__dlxtp_1
X_2225_ VGND VDPWR VDPWR VGND _0913_ _0791_ _1103_ _0786_ sky130_fd_sc_hd__mux2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[12\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[12\]\[1\] net237 dig_ctrl_inst.latch_mem_inst.gclk\[12\]
+ sky130_fd_sc_hd__dlxtp_1
Xclkbuf_leaf_18_clk VGND VDPWR VDPWR VGND clknet_leaf_18_clk clknet_1_0__leaf_clk
+ sky130_fd_sc_hd__clkbuf_8
X_2087_ VDPWR VGND VDPWR VGND _0779_ net157 _0778_ _0780_ sky130_fd_sc_hd__a21o_1
X_2156_ VDPWR VGND VDPWR VGND dig_ctrl_inst.cpu_inst.data\[2\] _0743_ _0847_ _0825_
+ net161 _0846_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_5_Right_5 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_54_338 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[5\].gen_latches\[3\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[5\]\[3\] net223 dig_ctrl_inst.latch_mem_inst.gclk\[5\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_26_Left_104 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2010_ VGND VDPWR VDPWR VGND _0278_ dig_ctrl_inst.latch_mem_inst.RAM\[5\]\[7\] _0690_
+ _0702_ _0708_ _0715_ sky130_fd_sc_hd__a2111o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[38\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[38\]\[6\] net195 dig_ctrl_inst.latch_mem_inst.gclk\[38\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_35_Left_113 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_44_Left_122 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[27\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[27\]\[4\] net212 dig_ctrl_inst.latch_mem_inst.gclk\[27\]
+ sky130_fd_sc_hd__dlxtp_1
X_1725_ VDPWR VGND VDPWR VGND _0427_ _0431_ _0429_ _0426_ _0435_ sky130_fd_sc_hd__or4_1
Xclkbuf_leaf_7_clk VGND VDPWR VDPWR VGND clknet_leaf_7_clk clknet_1_1__leaf_clk sky130_fd_sc_hd__clkbuf_8
Xhold103 VGND VDPWR VDPWR VGND net385 net19 sky130_fd_sc_hd__dlygate4sd3_1
X_1656_ VDPWR VGND VDPWR VGND _0367_ net64 net72 dig_ctrl_inst.latch_mem_inst.RAM\[30\]\[1\]
+ sky130_fd_sc_hd__and3_2
X_1587_ VGND VDPWR VDPWR VGND _0299_ net46 net81 net105 dig_ctrl_inst.latch_mem_inst.RAM\[63\]\[0\]
+ sky130_fd_sc_hd__and4_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[16\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[16\]\[2\] net225 dig_ctrl_inst.latch_mem_inst.gclk\[16\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_53_Left_131 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_28_91 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
X_2208_ VGND VDPWR VDPWR VGND _0787_ _0240_ _0786_ _1118_ _0897_ _0896_ sky130_fd_sc_hd__o221a_1
X_2139_ VGND VDPWR VDPWR VGND _0831_ _0748_ _0830_ _0750_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_187 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_62_Left_140 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[9\].gen_latches\[4\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[9\]\[4\] net212 dig_ctrl_inst.latch_mem_inst.gclk\[9\]
+ sky130_fd_sc_hd__dlxtp_1
X_2490_ VGND VDPWR VDPWR VGND clknet_leaf_5_clk _0089_ net178 dig_ctrl_inst.spi_data_i\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_1441_ VGND VDPWR VDPWR VGND net248 _1007_ dig_ctrl_inst.cpu_inst.prev_state\[2\]
+ _0999_ _0178_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_49_35 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
X_1510_ VDPWR VGND VDPWR VGND _0224_ _1005_ _1006_ _0216_ _0174_ _0223_ sky130_fd_sc_hd__o32a_1
X_1372_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[42\] net57 net83
+ net153 sky130_fd_sc_hd__and3_2
XFILLER_0_65_23 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_18_338 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[51\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[51\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[51\] sky130_fd_sc_hd__clkbuf_4
X_1708_ VDPWR VGND VDPWR VGND _0125_ dig_ctrl_inst.latch_mem_inst.RAM\[18\]\[2\] _0121_
+ _0418_ dig_ctrl_inst.latch_mem_inst.RAM\[22\]\[2\] sky130_fd_sc_hd__a22o_1
XFILLER_0_5_298 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
X_1639_ VDPWR VGND VDPWR VGND _0350_ net46 net96 dig_ctrl_inst.latch_mem_inst.RAM\[52\]\[1\]
+ sky130_fd_sc_hd__and3_2
Xfanout75 VGND VDPWR VDPWR VGND _0115_ net75 sky130_fd_sc_hd__clkbuf_2
Xfanout97 VDPWR VGND VDPWR VGND net97 net98 sky130_fd_sc_hd__buf_2
Xfanout42 VGND VDPWR VDPWR VGND net47 net42 sky130_fd_sc_hd__clkbuf_2
Xfanout86 VDPWR VGND VDPWR VGND net86 net87 sky130_fd_sc_hd__buf_2
Xfanout64 VDPWR VGND VDPWR VGND net64 net66 sky130_fd_sc_hd__buf_2
Xfanout53 VDPWR VGND VDPWR VGND net54 net53 sky130_fd_sc_hd__buf_4
XFILLER_0_51_149 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_51_69 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_27_113 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_1990_ VDPWR VGND VDPWR VGND _0695_ net61 net93 dig_ctrl_inst.latch_mem_inst.RAM\[22\]\[7\]
+ sky130_fd_sc_hd__and3_2
Xclkload12 VGND VDPWR VDPWR VGND clkload12/Y clknet_leaf_5_clk sky130_fd_sc_hd__inv_8
Xdig_ctrl_inst.latch_mem_inst.gen_words\[60\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[60\]\[4\] net209 dig_ctrl_inst.latch_mem_inst.gclk\[60\]
+ sky130_fd_sc_hd__dlxtp_1
X_2473_ VGND VDPWR VDPWR VGND clknet_leaf_4_clk _0079_ net174 dig_ctrl_inst.spi_data_o\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_193 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1355_ VDPWR VGND VDPWR VGND _0135_ net55 net116 net131 sky130_fd_sc_hd__and3_2
X_1424_ VDPWR VGND VDPWR VGND net255 dig_ctrl_inst.cpu_inst.r0\[6\] net259 _0166_
+ sky130_fd_sc_hd__or3_1
X_1286_ VDPWR VGND VDPWR VGND _1047_ net135 net134 net304 _1132_ _1078_ sky130_fd_sc_hd__a2111oi_1
Xclkload6 VDPWR VGND VDPWR VGND clkload6/Y clknet_leaf_16_clk sky130_fd_sc_hd__inv_6
Xfanout221 VDPWR VGND VDPWR VGND net221 net223 sky130_fd_sc_hd__dlymetal6s2s_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[12\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[12\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[12\] clknet_leaf_0_clk sky130_fd_sc_hd__dlclkp_1
X_2521__279 VGND VDPWR VDPWR VGND _2521__279/LO net279 sky130_fd_sc_hd__conb_1
Xfanout243 VGND VDPWR VDPWR VGND net244 net243 sky130_fd_sc_hd__clkbuf_2
Xfanout265 VDPWR VGND VDPWR VGND net266 net265 sky130_fd_sc_hd__buf_4
Xfanout254 VDPWR VGND VDPWR VGND net255 net254 sky130_fd_sc_hd__buf_4
Xfanout232 VGND VDPWR VDPWR VGND net233 net232 sky130_fd_sc_hd__clkbuf_2
Xfanout210 VGND VDPWR VDPWR VGND net323 net210 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_46_47 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_27 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_1973_ VDPWR VGND VDPWR VGND _0678_ _0677_ _0676_ _0675_ _0679_ sky130_fd_sc_hd__or4_4
X_2525_ VDPWR VGND VDPWR VGND uio_oe[6] net280 sky130_fd_sc_hd__buf_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[53\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[53\]\[3\] net216 dig_ctrl_inst.latch_mem_inst.gclk\[53\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_39_3 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_2387_ VGND VDPWR VDPWR VGND clknet_leaf_4_clk net330 net175 dig_ctrl_inst.synchronizer_port_i_inst\[3\].out
+ sky130_fd_sc_hd__dfrtp_1
X_2456_ VGND VDPWR VDPWR VGND clknet_leaf_6_clk _0064_ net145 dig_ctrl_inst.cpu_inst.r2\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_1338_ VDPWR VGND VDPWR VGND _0127_ net86 net64 sky130_fd_sc_hd__and2_1
X_1407_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[61\] net150 _0158_
+ sky130_fd_sc_hd__and2_1
X_1269_ VDPWR VGND VDPWR VGND net256 dig_ctrl_inst.cpu_inst.r0\[4\] net260 _1117_
+ sky130_fd_sc_hd__or3_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[42\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[42\]\[1\] net237 dig_ctrl_inst.latch_mem_inst.gclk\[42\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[44\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[44\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[44\] sky130_fd_sc_hd__clkbuf_4
X_2172_ VGND VDPWR VDPWR VGND _0768_ _0817_ net167 _0862_ sky130_fd_sc_hd__o21a_1
X_2241_ VGND VDPWR VDPWR VGND _0927_ _0230_ _0928_ sky130_fd_sc_hd__xnor2_1
X_2310_ VGND VDPWR VDPWR VGND _0070_ _0969_ _0977_ net358 sky130_fd_sc_hd__mux2_1
X_1956_ VGND VDPWR VDPWR VGND _0662_ net57 net73 dig_ctrl_inst.latch_mem_inst.RAM\[46\]\[6\]
+ _0145_ dig_ctrl_inst.latch_mem_inst.RAM\[45\]\[6\] sky130_fd_sc_hd__a32o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[57\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[57\]\[4\] net210 dig_ctrl_inst.latch_mem_inst.gclk\[57\]
+ sky130_fd_sc_hd__dlxtp_1
X_1887_ VDPWR VGND VDPWR VGND _0150_ dig_ctrl_inst.latch_mem_inst.RAM\[13\]\[5\] _0114_
+ _0594_ dig_ctrl_inst.latch_mem_inst.RAM\[52\]\[5\] sky130_fd_sc_hd__a22o_1
Xoutput19 VDPWR VGND VDPWR VGND port_ms_o[2] net19 sky130_fd_sc_hd__buf_2
X_2508_ VGND VDPWR VDPWR VGND clknet_leaf_5_clk _0105_ net178 net19 sky130_fd_sc_hd__dfrtp_1
X_2439_ VGND VDPWR VDPWR VGND clknet_leaf_8_clk _0047_ net146 dig_ctrl_inst.cpu_inst.r0\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[46\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[46\]\[2\] net228 dig_ctrl_inst.latch_mem_inst.gclk\[46\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[1\].gen_latches\[6\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[1\]\[6\] net195 dig_ctrl_inst.latch_mem_inst.gclk\[1\]
+ sky130_fd_sc_hd__dlxtp_1
X_2527__274 VGND VDPWR VDPWR VGND net274 _2527__274/HI sky130_fd_sc_hd__conb_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[35\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[35\]\[0\] net240 dig_ctrl_inst.latch_mem_inst.gclk\[35\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_43_15 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_1741_ VDPWR VGND VDPWR VGND _0146_ dig_ctrl_inst.latch_mem_inst.RAM\[44\]\[3\] _0144_
+ _0450_ dig_ctrl_inst.latch_mem_inst.RAM\[47\]\[3\] sky130_fd_sc_hd__a22o_1
X_1810_ VDPWR VGND VDPWR VGND _0513_ _0517_ _0512_ _0518_ sky130_fd_sc_hd__or3_1
X_1672_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[11\]\[1\] _1145_ _0383_
+ _0126_ dig_ctrl_inst.latch_mem_inst.RAM\[23\]\[1\] _0377_ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_333 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[23\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[23\]\[7\] net183 dig_ctrl_inst.latch_mem_inst.gclk\[23\]
+ sky130_fd_sc_hd__dlxtp_1
X_2224_ VGND VDPWR VDPWR VGND _0890_ net160 _0912_ sky130_fd_sc_hd__xnor2_1
X_2155_ VGND VDPWR VDPWR VGND _0783_ net169 _0786_ net168 _0846_ sky130_fd_sc_hd__a2bb2o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[12\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[12\]\[5\] net200 dig_ctrl_inst.latch_mem_inst.gclk\[12\]
+ sky130_fd_sc_hd__dlxtp_1
X_2086_ VGND VDPWR VDPWR VGND _0233_ _0779_ net137 sky130_fd_sc_hd__nand2_1
X_1939_ VDPWR VGND VDPWR VGND _0645_ net65 net84 dig_ctrl_inst.latch_mem_inst.RAM\[26\]\[6\]
+ sky130_fd_sc_hd__and3_2
XFILLER_0_16_244 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_31_225 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[5\].gen_latches\[7\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[5\]\[7\] net187 dig_ctrl_inst.latch_mem_inst.gclk\[5\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[39\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[39\]\[1\] net232 dig_ctrl_inst.latch_mem_inst.gclk\[39\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_11_Right_11 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[1\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[1\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[1\] sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_20_Right_20 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_60_309 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xhold104 VGND VDPWR VDPWR VGND net386 net20 sky130_fd_sc_hd__dlygate4sd3_1
X_1724_ VDPWR VGND VDPWR VGND _0419_ _0433_ _0423_ _0417_ _0434_ sky130_fd_sc_hd__or4_1
X_1586_ VDPWR VGND VDPWR VGND _0298_ net294 net121 dig_ctrl_inst.latch_mem_inst.RAM\[10\]\[0\]
+ sky130_fd_sc_hd__and3_2
X_1655_ VDPWR VGND VDPWR VGND _0366_ net61 net128 dig_ctrl_inst.latch_mem_inst.RAM\[16\]\[1\]
+ sky130_fd_sc_hd__and3_2
X_2138_ VDPWR VGND VDPWR VGND _0830_ _0828_ _0829_ sky130_fd_sc_hd__and2_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[17\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[17\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[17\] clknet_leaf_1_clk sky130_fd_sc_hd__dlclkp_1
XFILLER_0_48_111 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_3 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_81 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2069_ VGND VDPWR VDPWR VGND net166 _0762_ net137 sky130_fd_sc_hd__nand2_1
X_2207_ VDPWR VGND VDPWR VGND net169 _0825_ _0896_ _1118_ _0790_ sky130_fd_sc_hd__a22oi_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[16\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[16\]\[6\] net191 dig_ctrl_inst.latch_mem_inst.gclk\[16\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_63_125 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
X_1440_ VDPWR VGND VDPWR VGND dig_ctrl_inst.cpu_inst.prev_state\[2\] net248 _1007_
+ _0177_ _0999_ sky130_fd_sc_hd__a22o_1
X_1371_ VDPWR VGND VDPWR VGND net83 net60 _0142_ sky130_fd_sc_hd__and2_2
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[37\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[37\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[37\] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_45_136 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_69_3 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1638_ VDPWR VGND VDPWR VGND _0349_ net61 net109 dig_ctrl_inst.latch_mem_inst.RAM\[18\]\[1\]
+ sky130_fd_sc_hd__and3_2
X_1707_ VDPWR VGND VDPWR VGND _0136_ dig_ctrl_inst.latch_mem_inst.RAM\[24\]\[2\] _0127_
+ _0417_ dig_ctrl_inst.latch_mem_inst.RAM\[34\]\[2\] sky130_fd_sc_hd__a22o_1
X_1569_ VGND VDPWR VDPWR VGND _0281_ net108 _1048_ net123 sky130_fd_sc_hd__a21bo_1
XPHY_EDGE_ROW_18_Left_96 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xfanout98 VGND VDPWR VDPWR VGND _1137_ net98 sky130_fd_sc_hd__clkbuf_2
Xfanout65 VDPWR VGND VDPWR VGND net65 net66 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout54 VDPWR VGND VDPWR VGND net60 net54 sky130_fd_sc_hd__buf_6
Xfanout76 VGND VDPWR VDPWR VGND net79 net76 sky130_fd_sc_hd__clkbuf_2
Xfanout43 VGND VDPWR VDPWR VGND net44 net43 sky130_fd_sc_hd__clkbuf_2
Xfanout87 VDPWR VGND VDPWR VGND net87 _1141_ sky130_fd_sc_hd__buf_2
XFILLER_0_19_17 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_27_125 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
Xclkload13 VGND VDPWR VDPWR VGND clknet_leaf_6_clk clkload13/Y sky130_fd_sc_hd__clkinv_8
X_2472_ VDPWR VGND VDPWR VGND clknet_leaf_4_clk _0078_ dig_ctrl_inst.spi_receiver_inst.stb_o
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_180 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
X_1354_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[32\] net55 net150
+ net128 sky130_fd_sc_hd__and3_2
X_1285_ VDPWR VGND VDPWR VGND _1078_ net304 net301 _1131_ sky130_fd_sc_hd__a21oi_1
X_1423_ VGND VDPWR VDPWR VGND net255 _0165_ dig_ctrl_inst.cpu_inst.r1\[6\] sky130_fd_sc_hd__and2b_1
Xclkload7 VGND VDPWR VDPWR VGND clkload7/Y clknet_leaf_18_clk sky130_fd_sc_hd__inv_16
XFILLER_0_14_331 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_41_172 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
Xfanout222 VDPWR VGND VDPWR VGND net222 net223 sky130_fd_sc_hd__buf_2
Xfanout211 VGND VDPWR VDPWR VGND net213 net211 sky130_fd_sc_hd__clkbuf_2
Xfanout200 VDPWR VGND VDPWR VGND net200 net201 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout244 VGND VDPWR VDPWR VGND net245 net244 sky130_fd_sc_hd__clkbuf_2
Xfanout233 VGND VDPWR VDPWR VGND net327 net233 sky130_fd_sc_hd__clkbuf_2
Xfanout255 VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.arg1\[1\] net255 sky130_fd_sc_hd__clkbuf_2
Xfanout266 VDPWR VGND VDPWR VGND net266 dig_ctrl_inst.cpu_inst.arg0\[0\] sky130_fd_sc_hd__buf_2
XFILLER_0_46_59 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_1_39 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1972_ VGND VDPWR VDPWR VGND _0117_ dig_ctrl_inst.latch_mem_inst.RAM\[15\]\[6\] _0625_
+ _0636_ _0658_ _0678_ sky130_fd_sc_hd__a2111o_1
X_2455_ VGND VDPWR VDPWR VGND clknet_leaf_8_clk _0063_ net143 dig_ctrl_inst.cpu_inst.r2\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_49_Right_49 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2524_ VDPWR VGND VDPWR VGND uio_oe[5] net273 sky130_fd_sc_hd__buf_2
XFILLER_0_11_73 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_58_Right_58 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2386_ VGND VDPWR VDPWR VGND clknet_leaf_3_clk net6 net174 dig_ctrl_inst.synchronizer_port_i_inst\[3\].pipe\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_1268_ VGND VDPWR VDPWR VGND net256 _1116_ dig_ctrl_inst.cpu_inst.r1\[4\] sky130_fd_sc_hd__and2b_1
X_1337_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[23\] net150 _0126_
+ sky130_fd_sc_hd__and2_1
X_1406_ VDPWR VGND VDPWR VGND _0158_ net44 net80 net115 sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[53\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[53\]\[7\] net184 dig_ctrl_inst.latch_mem_inst.gclk\[53\]
+ sky130_fd_sc_hd__dlxtp_1
X_1199_ VGND VDPWR VDPWR VGND _1047_ _1008_ _1046_ _1038_ _1029_ net249 sky130_fd_sc_hd__o41a_4
XFILLER_0_14_172 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_67_Right_67 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[42\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[42\]\[5\] net205 dig_ctrl_inst.latch_mem_inst.gclk\[42\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_76_Right_76 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[31\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[31\]\[3\] net215 dig_ctrl_inst.latch_mem_inst.gclk\[31\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[20\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[20\]\[1\] net235 dig_ctrl_inst.latch_mem_inst.gclk\[20\]
+ sky130_fd_sc_hd__dlxtp_1
X_2171_ VGND VDPWR VDPWR VGND _0765_ _0808_ _0768_ _0816_ _0861_ sky130_fd_sc_hd__o22a_1
X_2240_ VDPWR VGND VDPWR VGND _0906_ _0244_ _0241_ _0927_ sky130_fd_sc_hd__a21oi_1
X_1955_ VDPWR VGND VDPWR VGND _0277_ dig_ctrl_inst.latch_mem_inst.RAM\[21\]\[6\] _0124_
+ _0661_ dig_ctrl_inst.latch_mem_inst.RAM\[4\]\[6\] sky130_fd_sc_hd__a22o_1
X_1886_ VDPWR VGND VDPWR VGND _0586_ _0592_ _0588_ _0582_ _0593_ sky130_fd_sc_hd__or4_1
XFILLER_0_7_147 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2507_ VGND VDPWR VDPWR VGND clknet_leaf_4_clk _0104_ net178 net18 sky130_fd_sc_hd__dfrtp_1
X_2438_ VGND VDPWR VDPWR VGND clknet_leaf_7_clk _0046_ net144 dig_ctrl_inst.cpu_inst.r0\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_2369_ VGND VDPWR VDPWR VGND _0996_ net252 _0175_ _1013_ net253 sky130_fd_sc_hd__and4b_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[2\].gen_latches\[1\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[2\]\[1\] net232 dig_ctrl_inst.latch_mem_inst.gclk\[2\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[46\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[46\]\[6\] net197 dig_ctrl_inst.latch_mem_inst.gclk\[46\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_6_191 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[35\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[35\]\[4\] net210 dig_ctrl_inst.latch_mem_inst.gclk\[35\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[24\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[24\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[24\] clknet_leaf_17_clk sky130_fd_sc_hd__dlclkp_1
XFILLER_0_57_337 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_43_27 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_43_49 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
Xdig_ctrl_inst.latch_mem_inst.gen_words\[24\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[24\]\[2\] net227 dig_ctrl_inst.latch_mem_inst.gclk\[24\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_6_Left_84 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1740_ VGND VDPWR VDPWR VGND _0028_ _0449_ _0276_ net261 sky130_fd_sc_hd__mux2_1
X_1671_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[3\]\[1\] _1135_ _0382_
+ _0130_ dig_ctrl_inst.latch_mem_inst.RAM\[27\]\[1\] _0378_ sky130_fd_sc_hd__a221o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[13\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[13\]\[0\] net246 dig_ctrl_inst.latch_mem_inst.gclk\[13\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_68_24 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2085_ VDPWR VGND VDPWR VGND net137 net138 net157 _0778_ sky130_fd_sc_hd__a21oi_1
X_2154_ VGND VDPWR VDPWR VGND _0845_ _0750_ _0844_ _0748_ sky130_fd_sc_hd__mux2_1
X_2223_ VDPWR VGND VDPWR VGND net159 _0867_ net160 _0911_ sky130_fd_sc_hd__or3_1
XFILLER_0_16_223 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_1938_ VDPWR VGND VDPWR VGND _0644_ net48 net88 dig_ctrl_inst.latch_mem_inst.RAM\[56\]\[6\]
+ sky130_fd_sc_hd__and3_2
X_1869_ VDPWR VGND VDPWR VGND _0277_ dig_ctrl_inst.latch_mem_inst.RAM\[29\]\[5\] _0131_
+ _0576_ dig_ctrl_inst.latch_mem_inst.RAM\[4\]\[5\] sky130_fd_sc_hd__a22o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[6\].gen_latches\[2\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[6\]\[2\] net226 dig_ctrl_inst.latch_mem_inst.gclk\[6\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_39_337 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[39\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[39\]\[5\] net206 dig_ctrl_inst.latch_mem_inst.gclk\[39\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[28\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[28\]\[3\] net222 dig_ctrl_inst.latch_mem_inst.gclk\[28\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[17\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[17\]\[1\] net239 dig_ctrl_inst.latch_mem_inst.gclk\[17\]
+ sky130_fd_sc_hd__dlxtp_1
X_1723_ VGND VDPWR VDPWR VGND _0433_ net58 net96 dig_ctrl_inst.latch_mem_inst.RAM\[36\]\[2\]
+ _0279_ dig_ctrl_inst.latch_mem_inst.RAM\[6\]\[2\] sky130_fd_sc_hd__a32o_1
X_1654_ VDPWR VGND VDPWR VGND _0365_ net294 net121 dig_ctrl_inst.latch_mem_inst.RAM\[10\]\[1\]
+ sky130_fd_sc_hd__and3_2
Xhold105 VGND VDPWR VDPWR VGND net387 dig_ctrl_inst.cpu_inst.data\[7\] sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_248 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_2206_ VDPWR VGND VDPWR VGND _0792_ _0238_ _0894_ _0895_ sky130_fd_sc_hd__a21oi_1
X_1585_ VGND VDPWR VDPWR VGND _0297_ net63 net90 net116 dig_ctrl_inst.latch_mem_inst.RAM\[25\]\[0\]
+ sky130_fd_sc_hd__and4_1
X_2137_ VGND VDPWR VDPWR VGND net165 _0829_ net162 sky130_fd_sc_hd__nand2_1
XFILLER_0_44_81 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2068_ VGND VDPWR VDPWR VGND net169 _0761_ net137 sky130_fd_sc_hd__nand2_1
XFILLER_0_14_3 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_39_189 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_24_29 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_49_48 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_1370_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[41\] net152 _0141_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_45_126 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_14_62 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1706_ VGND VDPWR VDPWR VGND _0416_ net101 net106 net126 dig_ctrl_inst.latch_mem_inst.RAM\[7\]\[2\]
+ sky130_fd_sc_hd__and4_1
X_1637_ VDPWR VGND VDPWR VGND _0348_ net54 net94 dig_ctrl_inst.latch_mem_inst.RAM\[38\]\[1\]
+ sky130_fd_sc_hd__and3_2
XFILLER_0_5_256 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
X_1568_ VGND VDPWR VDPWR VGND _0280_ net119 _1131_ net101 net123 sky130_fd_sc_hd__o211a_1
X_1499_ VGND VDPWR VDPWR VGND _0215_ dig_ctrl_inst.cpu_inst.ip\[3\] dig_ctrl_inst.cpu_inst.ip\[2\]
+ dig_ctrl_inst.cpu_inst.ip\[1\] dig_ctrl_inst.cpu_inst.ip\[0\] sky130_fd_sc_hd__and4_1
Xfanout55 VGND VDPWR VDPWR VGND net60 net55 sky130_fd_sc_hd__clkbuf_2
Xfanout44 VDPWR VGND VDPWR VGND net44 net47 sky130_fd_sc_hd__buf_2
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[3\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[3\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[3\] clknet_leaf_3_clk sky130_fd_sc_hd__dlclkp_1
Xfanout88 VDPWR VGND VDPWR VGND net88 net89 sky130_fd_sc_hd__buf_2
Xfanout77 VGND VDPWR VDPWR VGND net77 net79 sky130_fd_sc_hd__buf_1
Xfanout99 VGND VDPWR VDPWR VGND net100 net99 sky130_fd_sc_hd__clkbuf_4
Xfanout66 VDPWR VGND VDPWR VGND net67 net66 sky130_fd_sc_hd__buf_4
XFILLER_0_3_3 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
Xdig_ctrl_inst.latch_mem_inst.gen_words\[61\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[61\]\[3\] net215 dig_ctrl_inst.latch_mem_inst.gclk\[61\]
+ sky130_fd_sc_hd__dlxtp_1
X_2471_ VGND VDPWR VDPWR VGND clknet_leaf_3_clk _0077_ net173 dig_ctrl_inst.spi_miso_o
+ sky130_fd_sc_hd__dfrtp_1
Xclkload14 VGND VDPWR VDPWR VGND clkload14/Y clknet_leaf_7_clk sky130_fd_sc_hd__clkinv_16
XFILLER_0_23_332 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1422_ VGND VDPWR VDPWR VGND net259 _0164_ dig_ctrl_inst.cpu_inst.r2\[6\] sky130_fd_sc_hd__and2b_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[50\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[50\]\[1\] net232 dig_ctrl_inst.latch_mem_inst.gclk\[50\]
+ sky130_fd_sc_hd__dlxtp_1
X_1284_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[1\] net154 _1130_
+ sky130_fd_sc_hd__and2_1
X_1353_ VDPWR VGND VDPWR VGND net129 net53 _0134_ sky130_fd_sc_hd__and2_2
Xclkload8 VGND VDPWR VDPWR VGND clkload8/Y clknet_leaf_1_clk sky130_fd_sc_hd__inv_12
XFILLER_0_41_71 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xfanout212 VGND VDPWR VDPWR VGND net213 net212 sky130_fd_sc_hd__clkbuf_2
Xfanout223 VDPWR VGND VDPWR VGND net223 net329 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout256 VDPWR VGND VDPWR VGND net257 net256 sky130_fd_sc_hd__buf_4
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[29\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[29\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[29\] clknet_leaf_0_clk sky130_fd_sc_hd__dlclkp_1
Xfanout245 VGND VDPWR VDPWR VGND net246 net245 sky130_fd_sc_hd__clkbuf_2
Xfanout234 VGND VDPWR VDPWR VGND net236 net234 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_1_281 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
Xfanout201 VGND VDPWR VDPWR VGND net202 net201 sky130_fd_sc_hd__clkbuf_2
Xfanout267 VDPWR VGND VDPWR VGND net268 net267 sky130_fd_sc_hd__buf_4
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[31\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[31\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[31\] clknet_leaf_15_clk sky130_fd_sc_hd__dlclkp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[54\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[54\]\[2\] net224 dig_ctrl_inst.latch_mem_inst.gclk\[54\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_23_140 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1971_ VGND VDPWR VDPWR VGND _0114_ dig_ctrl_inst.latch_mem_inst.RAM\[13\]\[6\] _0630_
+ _0641_ _0657_ _0677_ sky130_fd_sc_hd__a2111o_1
X_2385_ VGND VDPWR VDPWR VGND clknet_leaf_4_clk net332 net174 dig_ctrl_inst.synchronizer_port_i_inst\[4\].out
+ sky130_fd_sc_hd__dfrtp_1
X_2520__270 VGND VDPWR VDPWR VGND net270 _2520__270/HI sky130_fd_sc_hd__conb_1
X_2523_ VDPWR VGND VDPWR VGND uio_oe[4] net272 sky130_fd_sc_hd__buf_2
X_1405_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[60\] net48 net78
+ net153 sky130_fd_sc_hd__and3_2
X_2454_ VGND VDPWR VDPWR VGND clknet_leaf_9_clk _0062_ net141 dig_ctrl_inst.cpu_inst.r2\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_1336_ VGND VDPWR VDPWR VGND _0126_ net102 net99 net63 sky130_fd_sc_hd__and3_4
X_1267_ VGND VDPWR VDPWR VGND net256 net260 _1115_ dig_ctrl_inst.cpu_inst.r2\[4\]
+ sky130_fd_sc_hd__and3b_1
X_1198_ VDPWR VGND VDPWR VGND _1046_ _1039_ _1045_ sky130_fd_sc_hd__and2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[43\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[43\]\[0\] net245 dig_ctrl_inst.latch_mem_inst.gclk\[43\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_36_71 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xinput1 VGND VDPWR VDPWR VGND net1 port_ms_i sky130_fd_sc_hd__buf_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[31\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[31\]\[7\] net187 dig_ctrl_inst.latch_mem_inst.gclk\[31\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_32_29 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[20\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[20\]\[5\] net207 dig_ctrl_inst.latch_mem_inst.gclk\[20\]
+ sky130_fd_sc_hd__dlxtp_1
X_2170_ VGND VDPWR VDPWR VGND _0770_ _0836_ _0809_ _0859_ _0860_ sky130_fd_sc_hd__o22a_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[58\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[58\]\[3\] net223 dig_ctrl_inst.latch_mem_inst.gclk\[58\]
+ sky130_fd_sc_hd__dlxtp_1
X_1954_ VDPWR VGND VDPWR VGND _0153_ dig_ctrl_inst.latch_mem_inst.RAM\[22\]\[6\] _0125_
+ _0660_ dig_ctrl_inst.latch_mem_inst.RAM\[55\]\[6\] sky130_fd_sc_hd__a22o_1
X_1885_ VGND VDPWR VDPWR VGND _1135_ dig_ctrl_inst.latch_mem_inst.RAM\[3\]\[5\] _0589_
+ _0590_ _0591_ _0592_ sky130_fd_sc_hd__a2111o_1
X_2506_ VGND VDPWR VDPWR VGND clknet_leaf_3_clk _0103_ net178 net17 sky130_fd_sc_hd__dfrtp_1
X_2437_ VGND VDPWR VDPWR VGND clknet_leaf_7_clk _0045_ net144 dig_ctrl_inst.cpu_inst.r0\[0\]
+ sky130_fd_sc_hd__dfrtp_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[47\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[47\]\[1\] net236 dig_ctrl_inst.latch_mem_inst.gclk\[47\]
+ sky130_fd_sc_hd__dlxtp_1
X_2368_ VGND VDPWR VDPWR VGND _0991_ _0566_ _0992_ _0993_ _0994_ _0995_ sky130_fd_sc_hd__a2111o_1
X_1319_ VGND VDPWR VDPWR VGND _0117_ net126 net106 net82 sky130_fd_sc_hd__and3_4
X_2299_ VGND VDPWR VDPWR VGND _0976_ _1024_ _0175_ _0756_ sky130_fd_sc_hd__and3_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[2\].gen_latches\[5\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[2\]\[5\] net203 dig_ctrl_inst.latch_mem_inst.gclk\[2\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_6_181 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xmax_cap85 VDPWR VGND VDPWR VGND net85 _1144_ sky130_fd_sc_hd__dlymetal6s2s_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[24\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[24\]\[6\] net194 dig_ctrl_inst.latch_mem_inst.gclk\[24\]
+ sky130_fd_sc_hd__dlxtp_1
X_1670_ VGND VDPWR VDPWR VGND _0153_ dig_ctrl_inst.latch_mem_inst.RAM\[55\]\[1\] _0341_
+ _0359_ _0360_ _0381_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_68_36 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2222_ VDPWR VGND VDPWR VGND net167 _0810_ _0910_ _0819_ _0909_ net171 sky130_fd_sc_hd__a221o_1
XFILLER_0_48_316 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[13\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[13\]\[4\] net211 dig_ctrl_inst.latch_mem_inst.gclk\[13\]
+ sky130_fd_sc_hd__dlxtp_1
X_2084_ VGND VDPWR VDPWR VGND _0777_ _0776_ _1068_ _0775_ sky130_fd_sc_hd__mux2_1
X_2153_ VGND VDPWR VDPWR VGND _0842_ _0844_ _0843_ sky130_fd_sc_hd__nand2_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[40\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[40\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[40\] sky130_fd_sc_hd__clkbuf_4
X_1937_ VDPWR VGND VDPWR VGND _0643_ net55 net110 dig_ctrl_inst.latch_mem_inst.RAM\[34\]\[6\]
+ sky130_fd_sc_hd__and3_2
X_1799_ VDPWR VGND VDPWR VGND _0127_ dig_ctrl_inst.latch_mem_inst.RAM\[17\]\[4\] _0120_
+ _0507_ dig_ctrl_inst.latch_mem_inst.RAM\[24\]\[4\] sky130_fd_sc_hd__a22o_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[8\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[8\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[8\] clknet_leaf_3_clk sky130_fd_sc_hd__dlclkp_1
X_1868_ VDPWR VGND VDPWR VGND _0279_ dig_ctrl_inst.latch_mem_inst.RAM\[59\]\[5\] _0156_
+ _0575_ dig_ctrl_inst.latch_mem_inst.RAM\[6\]\[5\] sky130_fd_sc_hd__a22o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[6\].gen_latches\[6\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[6\]\[6\] net194 dig_ctrl_inst.latch_mem_inst.gclk\[6\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_15_290 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[28\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[28\]\[7\] net185 dig_ctrl_inst.latch_mem_inst.gclk\[28\]
+ sky130_fd_sc_hd__dlxtp_1
X_1722_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[51\]\[2\] _0149_ _0432_
+ _0277_ dig_ctrl_inst.latch_mem_inst.RAM\[4\]\[2\] _0402_ sky130_fd_sc_hd__a221o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[17\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[17\]\[5\] net202 dig_ctrl_inst.latch_mem_inst.gclk\[17\]
+ sky130_fd_sc_hd__dlxtp_1
X_1584_ VDPWR VGND VDPWR VGND _0296_ net63 net76 dig_ctrl_inst.latch_mem_inst.RAM\[28\]\[0\]
+ sky130_fd_sc_hd__and3_2
X_1653_ VDPWR VGND VDPWR VGND _0364_ net56 net96 dig_ctrl_inst.latch_mem_inst.RAM\[36\]\[1\]
+ sky130_fd_sc_hd__and3_2
XPHY_EDGE_ROW_9_Right_9 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xhold106 VGND VDPWR VDPWR VGND net388 dig_ctrl_inst.cpu_inst.data\[6\] sky130_fd_sc_hd__dlygate4sd3_1
X_2205_ VDPWR VGND VDPWR VGND _0783_ dig_ctrl_inst.cpu_inst.data\[4\] _0743_ _0894_
+ net160 sky130_fd_sc_hd__a22o_1
X_2136_ VGND VDPWR VDPWR VGND _0828_ net165 net162 sky130_fd_sc_hd__or2_1
XFILLER_0_48_135 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_48_168 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_22_Left_100 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_8_210 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2067_ VDPWR VGND VDPWR VGND _1118_ _0172_ _0167_ _1103_ _0760_ sky130_fd_sc_hd__or4_2
XFILLER_0_39_113 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[36\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[36\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[36\] clknet_leaf_19_clk sky130_fd_sc_hd__dlclkp_1
X_1705_ VDPWR VGND VDPWR VGND _0415_ net54 net77 dig_ctrl_inst.latch_mem_inst.RAM\[44\]\[2\]
+ sky130_fd_sc_hd__and3_2
X_1636_ VDPWR VGND VDPWR VGND _0347_ net46 net130 dig_ctrl_inst.latch_mem_inst.RAM\[48\]\[1\]
+ sky130_fd_sc_hd__and3_2
X_1567_ VDPWR VGND VDPWR VGND net125 net95 _0279_ sky130_fd_sc_hd__and2_2
X_2119_ VGND VDPWR VDPWR VGND _0811_ _0766_ _1068_ _0762_ sky130_fd_sc_hd__mux2_1
X_1498_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.ip\[2\] _0211_ _0204_ _0214_
+ _0021_ sky130_fd_sc_hd__a2bb2o_1
Xfanout78 VDPWR VGND VDPWR VGND net78 net79 sky130_fd_sc_hd__buf_2
Xfanout45 VDPWR VGND VDPWR VGND net45 net47 sky130_fd_sc_hd__buf_2
Xfanout67 VDPWR VGND VDPWR VGND _0118_ net67 sky130_fd_sc_hd__buf_4
Xfanout56 VGND VDPWR VDPWR VGND net60 net56 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_44_160 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
Xclkload15 VGND VDPWR VDPWR VGND clkload15/Y clknet_leaf_8_clk sky130_fd_sc_hd__inv_12
Xdig_ctrl_inst.latch_mem_inst.gen_words\[61\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[61\]\[7\] net184 dig_ctrl_inst.latch_mem_inst.gclk\[61\]
+ sky130_fd_sc_hd__dlxtp_1
X_2470_ VGND VDPWR VDPWR VGND clknet_leaf_11_clk _0076_ net140 dig_ctrl_inst.cpu_inst.r3\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_1421_ VDPWR VGND VDPWR VGND _0163_ dig_ctrl_inst.cpu_inst.r3\[6\] net255 net259
+ sky130_fd_sc_hd__and3_2
X_1352_ VGND VDPWR VDPWR VGND _1127_ _0133_ _1112_ sky130_fd_sc_hd__and2b_1
X_1283_ VDPWR VGND VDPWR VGND _1130_ net118 net125 net132 sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[50\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[50\]\[5\] net203 dig_ctrl_inst.latch_mem_inst.gclk\[50\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[33\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[33\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[33\] sky130_fd_sc_hd__clkbuf_4
Xclkload9 VGND VDPWR VDPWR VGND clkload9/Y clknet_leaf_2_clk sky130_fd_sc_hd__inv_16
Xfanout202 VDPWR VGND VDPWR VGND net202 net207 sky130_fd_sc_hd__buf_2
Xfanout257 VDPWR VGND VDPWR VGND net257 dig_ctrl_inst.cpu_inst.arg1\[1\] sky130_fd_sc_hd__buf_2
Xfanout246 VDPWR VGND VDPWR VGND net246 net247 sky130_fd_sc_hd__buf_2
Xfanout213 VDPWR VGND VDPWR VGND net213 net214 sky130_fd_sc_hd__buf_2
Xfanout268 VDPWR VGND VDPWR VGND dig_ctrl_inst.cpu_inst.arg0\[0\] net268 sky130_fd_sc_hd__buf_4
X_1619_ VDPWR VGND VDPWR VGND _0328_ _0330_ _0329_ _0327_ _0331_ sky130_fd_sc_hd__or4_1
Xfanout224 VGND VDPWR VDPWR VGND net225 net224 sky130_fd_sc_hd__clkbuf_2
Xfanout235 VGND VDPWR VDPWR VGND net235 net236 sky130_fd_sc_hd__buf_1
X_1970_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[31\]\[6\] _0132_ _0676_
+ _0134_ dig_ctrl_inst.latch_mem_inst.RAM\[32\]\[6\] _0643_ sky130_fd_sc_hd__a221o_1
X_2522_ VDPWR VGND VDPWR VGND uio_oe[3] net271 sky130_fd_sc_hd__buf_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[54\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[54\]\[6\] net191 dig_ctrl_inst.latch_mem_inst.gclk\[54\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_15_119 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_2384_ VGND VDPWR VDPWR VGND clknet_leaf_3_clk net7 net174 dig_ctrl_inst.synchronizer_port_i_inst\[4\].pipe\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_1404_ VDPWR VGND VDPWR VGND net78 net49 _0157_ sky130_fd_sc_hd__and2_2
X_1335_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[22\] net61 net93
+ net149 sky130_fd_sc_hd__and3_2
X_2453_ VGND VDPWR VDPWR VGND clknet_leaf_11_clk _0061_ net140 dig_ctrl_inst.cpu_inst.r2\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[43\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[43\]\[4\] net213 dig_ctrl_inst.latch_mem_inst.gclk\[43\]
+ sky130_fd_sc_hd__dlxtp_1
Xinput2 VGND VDPWR VDPWR VGND net2 rst_n sky130_fd_sc_hd__clkbuf_1
X_1266_ VDPWR VGND VDPWR VGND _1114_ dig_ctrl_inst.cpu_inst.r3\[4\] net256 net261
+ sky130_fd_sc_hd__and3_2
X_1197_ VGND VDPWR VDPWR VGND net300 _1041_ _1042_ _1043_ _1044_ _1045_ sky130_fd_sc_hd__o41a_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[32\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[32\]\[2\] net224 dig_ctrl_inst.latch_mem_inst.gclk\[32\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[21\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[21\]\[0\] net246 dig_ctrl_inst.latch_mem_inst.gclk\[21\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_69_Left_147 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[58\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[58\]\[7\] net188 dig_ctrl_inst.latch_mem_inst.gclk\[58\]
+ sky130_fd_sc_hd__dlxtp_1
X_1953_ VDPWR VGND VDPWR VGND _0659_ net50 net73 dig_ctrl_inst.latch_mem_inst.RAM\[62\]\[6\]
+ sky130_fd_sc_hd__and3_2
XFILLER_0_22_85 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1884_ VDPWR VGND VDPWR VGND _0591_ net44 net128 dig_ctrl_inst.latch_mem_inst.RAM\[48\]\[5\]
+ sky130_fd_sc_hd__and3_2
X_2505_ VGND VDPWR VDPWR VGND clknet_leaf_5_clk _0102_ net178 net35 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_333 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2436_ VDPWR VGND VDPWR VGND clknet_leaf_9_clk _0044_ dig_ctrl_inst.cpu_inst.prev_state\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[3\].gen_latches\[0\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[3\]\[0\] net243 dig_ctrl_inst.latch_mem_inst.gclk\[3\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_47_93 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
Xdig_ctrl_inst.latch_mem_inst.gen_words\[47\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[47\]\[5\] net203 dig_ctrl_inst.latch_mem_inst.gclk\[47\]
+ sky130_fd_sc_hd__dlxtp_1
X_2367_ VDPWR VGND VDPWR VGND _0994_ _0449_ _0623_ sky130_fd_sc_hd__and2_1
X_2298_ VGND VDPWR VDPWR VGND _0060_ _0975_ _0967_ net377 sky130_fd_sc_hd__mux2_1
X_1318_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[14\] net72 net120
+ net148 sky130_fd_sc_hd__and3_2
X_1249_ VGND VDPWR VDPWR VGND _1040_ _1097_ _1096_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_339 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[36\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[36\]\[3\] net218 dig_ctrl_inst.latch_mem_inst.gclk\[36\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_input_latches\[1\].n_latch VGND VDPWR VDPWR VGND
+ dig_ctrl_inst.latch_mem_inst.wdata\[1\] dig_ctrl_inst.data_out\[1\] clknet_leaf_2_clk
+ sky130_fd_sc_hd__dlxtn_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[25\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[25\]\[1\] net232 dig_ctrl_inst.latch_mem_inst.gclk\[25\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_25_225 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_68_15 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[43\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[43\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[43\] clknet_1_1__leaf_clk sky130_fd_sc_hd__dlclkp_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[26\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[26\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[26\] sky130_fd_sc_hd__clkbuf_4
X_2221_ VGND VDPWR VDPWR VGND _0908_ _0770_ _0859_ _0836_ _0909_ _0886_ sky130_fd_sc_hd__o221a_1
X_2152_ VGND VDPWR VDPWR VGND net161 net166 _0843_ net164 sky130_fd_sc_hd__o21ai_1
X_2083_ VGND VDPWR VDPWR VGND net159 _0776_ net137 sky130_fd_sc_hd__nand2_1
X_1867_ VGND VDPWR VDPWR VGND _1142_ dig_ctrl_inst.latch_mem_inst.RAM\[8\]\[5\] _0571_
+ _0572_ _0573_ _0574_ sky130_fd_sc_hd__a2111o_1
X_1936_ VDPWR VGND VDPWR VGND _0642_ net94 net121 dig_ctrl_inst.latch_mem_inst.RAM\[6\]\[6\]
+ sky130_fd_sc_hd__and3_2
X_1798_ VGND VDPWR VDPWR VGND _0029_ _0505_ _0276_ net257 sky130_fd_sc_hd__mux2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[7\].gen_latches\[1\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[7\]\[1\] net239 dig_ctrl_inst.latch_mem_inst.gclk\[7\]
+ sky130_fd_sc_hd__dlxtp_1
X_2419_ VGND VDPWR VDPWR VGND clknet_leaf_8_clk _0027_ net143 dig_ctrl_inst.cpu_inst.arg0\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_306 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_29 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[29\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[29\]\[2\] net229 dig_ctrl_inst.latch_mem_inst.gclk\[29\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[18\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[18\]\[0\] net242 dig_ctrl_inst.latch_mem_inst.gclk\[18\]
+ sky130_fd_sc_hd__dlxtp_1
X_1721_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[40\]\[2\] _0140_ _0431_
+ _0153_ dig_ctrl_inst.latch_mem_inst.RAM\[55\]\[2\] _0430_ sky130_fd_sc_hd__a221o_1
Xhold107 VGND VDPWR VDPWR VGND net389 net29 sky130_fd_sc_hd__dlygate4sd3_1
X_1583_ VGND VDPWR VDPWR VGND _0295_ net66 net91 net104 dig_ctrl_inst.latch_mem_inst.RAM\[27\]\[0\]
+ sky130_fd_sc_hd__and4_1
X_1652_ VDPWR VGND VDPWR VGND _0363_ net93 net120 dig_ctrl_inst.latch_mem_inst.RAM\[6\]\[1\]
+ sky130_fd_sc_hd__and3_2
X_2204_ VGND VDPWR VDPWR VGND _0747_ _0893_ _0892_ sky130_fd_sc_hd__nand2_1
X_2135_ VDPWR VGND VDPWR VGND _0783_ net166 _0826_ _0827_ sky130_fd_sc_hd__a21oi_1
X_2066_ VGND VDPWR VDPWR VGND _0759_ _0172_ _0167_ _1118_ _1103_ sky130_fd_sc_hd__nor4_1
X_1919_ VDPWR VGND VDPWR VGND _0625_ net44 net93 dig_ctrl_inst.latch_mem_inst.RAM\[54\]\[6\]
+ sky130_fd_sc_hd__and3_2
XFILLER_0_39_125 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1704_ VGND VDPWR VDPWR VGND _0414_ net69 _1146_ net119 dig_ctrl_inst.latch_mem_inst.RAM\[29\]\[2\]
+ sky130_fd_sc_hd__and4_1
XFILLER_0_30_85 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_5_214 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1566_ VDPWR VGND VDPWR VGND _0278_ net101 net118 net125 sky130_fd_sc_hd__and3_2
X_1497_ VDPWR VGND VDPWR VGND _0213_ _0173_ _0212_ _0214_ sky130_fd_sc_hd__a21oi_1
X_1635_ VDPWR VGND VDPWR VGND _0346_ net55 net109 dig_ctrl_inst.latch_mem_inst.RAM\[34\]\[1\]
+ sky130_fd_sc_hd__and3_2
X_2049_ VGND VDPWR VDPWR VGND net252 _0742_ net253 sky130_fd_sc_hd__nand2_1
X_2118_ VGND VDPWR VDPWR VGND _0810_ _0770_ _0809_ sky130_fd_sc_hd__or2_1
Xfanout68 VDPWR VGND VDPWR VGND net68 net71 sky130_fd_sc_hd__buf_2
Xfanout79 VDPWR VGND VDPWR VGND net79 _1147_ sky130_fd_sc_hd__buf_2
Xfanout57 VDPWR VGND VDPWR VGND net59 net57 sky130_fd_sc_hd__buf_4
Xfanout46 VGND VDPWR VDPWR VGND net47 net46 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_44_172 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
Xdig_ctrl_inst.latch_mem_inst.gen_words\[62\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[62\]\[2\] net230 dig_ctrl_inst.latch_mem_inst.gclk\[62\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_41_Left_119 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[51\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[51\]\[0\] net241 dig_ctrl_inst.latch_mem_inst.gclk\[51\]
+ sky130_fd_sc_hd__dlxtp_1
Xclkload16 VGND VDPWR VDPWR VGND clkload16/Y clknet_leaf_9_clk sky130_fd_sc_hd__inv_12
X_1420_ VDPWR VGND VDPWR VGND _1103_ net250 dig_ctrl_inst.spi_data_o\[5\] dig_ctrl_inst.data_out\[5\]
+ _0162_ sky130_fd_sc_hd__a22o_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[19\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[19\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[19\] sky130_fd_sc_hd__clkbuf_4
X_1351_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[31\] net151 _0132_
+ sky130_fd_sc_hd__and2_1
X_1282_ VGND VDPWR VDPWR VGND _1129_ _1076_ _1078_ net134 sky130_fd_sc_hd__and3_4
XPHY_EDGE_ROW_50_Left_128 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1618_ VDPWR VGND VDPWR VGND _0131_ dig_ctrl_inst.latch_mem_inst.RAM\[17\]\[0\] _0120_
+ _0330_ dig_ctrl_inst.latch_mem_inst.RAM\[29\]\[0\] sky130_fd_sc_hd__a22o_1
Xfanout247 VGND VDPWR VDPWR VGND net247 net325 sky130_fd_sc_hd__buf_1
Xfanout214 VDPWR VGND VDPWR VGND net214 net323 sky130_fd_sc_hd__buf_2
XFILLER_0_66_81 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xfanout203 VGND VDPWR VDPWR VGND net207 net203 sky130_fd_sc_hd__clkbuf_2
Xfanout236 VGND VDPWR VDPWR VGND net327 net236 sky130_fd_sc_hd__clkbuf_2
X_1549_ VDPWR VGND VDPWR VGND _0261_ _0253_ _0245_ _0262_ _0257_ sky130_fd_sc_hd__or4b_1
Xfanout225 VDPWR VGND VDPWR VGND net225 net231 sky130_fd_sc_hd__buf_2
Xfanout258 VDPWR VGND VDPWR VGND net259 net258 sky130_fd_sc_hd__buf_4
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[48\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[48\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[48\] clknet_leaf_12_clk sky130_fd_sc_hd__dlclkp_1
XFILLER_0_46_18 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
Xdig_ctrl_inst.latch_mem_inst.gen_words\[55\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[55\]\[1\] net233 dig_ctrl_inst.latch_mem_inst.gclk\[55\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_55_256 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_7_309 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
X_2521_ VDPWR VGND VDPWR VGND uio_oe[2] net279 sky130_fd_sc_hd__buf_2
XFILLER_0_11_337 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1265_ VGND VDPWR VDPWR VGND _1113_ net182 _1026_ _1027_ dig_ctrl_inst.cpu_inst.ip\[4\]
+ sky130_fd_sc_hd__o211a_1
X_2383_ VGND VDPWR VDPWR VGND clknet_leaf_4_clk net331 net174 dig_ctrl_inst.synchronizer_port_i_inst\[5\].out
+ sky130_fd_sc_hd__dfrtp_1
X_1403_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[59\] net153 _0156_
+ sky130_fd_sc_hd__and2_1
X_1334_ VDPWR VGND VDPWR VGND _0125_ net95 net68 sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_18_Right_18 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2452_ VGND VDPWR VDPWR VGND clknet_leaf_11_clk _0060_ net140 dig_ctrl_inst.cpu_inst.r1\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput3 VGND VDPWR VDPWR VGND net3 ui_in[0] sky130_fd_sc_hd__clkbuf_1
X_1196_ VDPWR VGND VDPWR VGND net264 dig_ctrl_inst.cpu_inst.r0\[3\] net268 _1044_
+ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_27_Right_27 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[50\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[50\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[50\] clknet_leaf_16_clk sky130_fd_sc_hd__dlclkp_1
XPHY_EDGE_ROW_36_Right_36 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[32\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[32\]\[6\] net191 dig_ctrl_inst.latch_mem_inst.gclk\[32\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_45_Right_45 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[21\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[21\]\[4\] net210 dig_ctrl_inst.latch_mem_inst.gclk\[21\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_54_Right_54 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[10\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[10\]\[2\] net228 dig_ctrl_inst.latch_mem_inst.gclk\[10\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[59\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[59\]\[2\] net230 dig_ctrl_inst.latch_mem_inst.gclk\[59\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_63_Right_63 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[48\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[48\]\[0\] net241 dig_ctrl_inst.latch_mem_inst.gclk\[48\]
+ sky130_fd_sc_hd__dlxtp_1
X_1952_ VGND VDPWR VDPWR VGND _0658_ net62 net100 net102 dig_ctrl_inst.latch_mem_inst.RAM\[23\]\[6\]
+ sky130_fd_sc_hd__and4_1
X_1883_ VDPWR VGND VDPWR VGND _0590_ net55 net75 dig_ctrl_inst.latch_mem_inst.RAM\[46\]\[5\]
+ sky130_fd_sc_hd__and3_2
X_2504_ VGND VDPWR VDPWR VGND clknet_leaf_5_clk _0101_ net178 net34 sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_72_Right_72 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2435_ VDPWR VGND VDPWR VGND clknet_leaf_8_clk _0043_ dig_ctrl_inst.cpu_inst.prev_state\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_2366_ VGND VDPWR VDPWR VGND _1009_ _0993_ _0685_ _0740_ sky130_fd_sc_hd__or3b_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[3\].gen_latches\[4\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[3\]\[4\] net212 dig_ctrl_inst.latch_mem_inst.gclk\[3\]
+ sky130_fd_sc_hd__dlxtp_1
X_1248_ VGND VDPWR VDPWR VGND net251 _1096_ dig_ctrl_inst.spi_receiver_inst.stb_o
+ sky130_fd_sc_hd__nand2_1
X_1317_ VDPWR VGND VDPWR VGND _0116_ net123 net73 sky130_fd_sc_hd__and2_1
XFILLER_0_2_41 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2297_ VGND VDPWR VDPWR VGND _0964_ _0963_ _0975_ _0751_ sky130_fd_sc_hd__o21ai_1
X_1179_ VGND VDPWR VDPWR VGND _1010_ net182 _1027_ sky130_fd_sc_hd__or2_4
XFILLER_0_63_82 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XANTENNA_30 VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_data_i\[0\] sky130_fd_sc_hd__diode_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[36\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[36\]\[7\] net185 dig_ctrl_inst.latch_mem_inst.gclk\[36\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[25\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[25\]\[5\] net203 dig_ctrl_inst.latch_mem_inst.gclk\[25\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_input_latches\[5\].n_latch VGND VDPWR VDPWR VGND
+ dig_ctrl_inst.latch_mem_inst.wdata\[5\] dig_ctrl_inst.data_out\[5\] clknet_leaf_8_clk
+ sky130_fd_sc_hd__dlxtn_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[14\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[14\]\[3\] net220 dig_ctrl_inst.latch_mem_inst.gclk\[14\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_0_337 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2220_ VGND VDPWR VDPWR VGND _0815_ _1068_ _0776_ _0908_ sky130_fd_sc_hd__o21ba_1
X_2151_ VDPWR VGND VDPWR VGND net164 net161 net166 _0842_ sky130_fd_sc_hd__or3_1
X_2082_ VGND VDPWR VDPWR VGND net160 _0775_ net137 sky130_fd_sc_hd__nand2_1
XFILLER_0_48_329 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1797_ VGND VDPWR VDPWR VGND net39 _0504_ _0288_ dig_ctrl_inst.latch_mem_inst.RAM\[0\]\[3\]
+ _0506_ sky130_fd_sc_hd__a2bb2o_1
X_1866_ VDPWR VGND VDPWR VGND _0573_ net59 net95 dig_ctrl_inst.latch_mem_inst.RAM\[38\]\[5\]
+ sky130_fd_sc_hd__and3_2
X_1935_ VGND VDPWR VDPWR VGND _0641_ net43 net90 net116 dig_ctrl_inst.latch_mem_inst.RAM\[57\]\[6\]
+ sky130_fd_sc_hd__and4_1
X_2418_ VGND VDPWR VDPWR VGND clknet_leaf_8_clk _0026_ net143 dig_ctrl_inst.cpu_inst.arg0\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_71 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[7\].gen_latches\[5\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[7\]\[5\] net206 dig_ctrl_inst.latch_mem_inst.gclk\[7\]
+ sky130_fd_sc_hd__dlxtp_1
X_2349_ VGND VDPWR VDPWR VGND _0099_ net32 _0987_ dig_ctrl_inst.cpu_inst.port_o\[4\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_318 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_0_Right_0 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_30_262 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[29\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[29\]\[6\] net197 dig_ctrl_inst.latch_mem_inst.gclk\[29\]
+ sky130_fd_sc_hd__dlxtp_1
Xhold108 VGND VDPWR VDPWR VGND net390 net28 sky130_fd_sc_hd__dlygate4sd3_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[18\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[18\]\[4\] net213 dig_ctrl_inst.latch_mem_inst.gclk\[18\]
+ sky130_fd_sc_hd__dlxtp_1
X_1720_ VDPWR VGND VDPWR VGND _0150_ dig_ctrl_inst.latch_mem_inst.RAM\[23\]\[2\] _0126_
+ _0430_ dig_ctrl_inst.latch_mem_inst.RAM\[52\]\[2\] sky130_fd_sc_hd__a22o_1
X_1651_ VDPWR VGND VDPWR VGND _0362_ net66 net294 dig_ctrl_inst.latch_mem_inst.RAM\[26\]\[1\]
+ sky130_fd_sc_hd__and3_2
X_1582_ VDPWR VGND VDPWR VGND _0294_ net48 net73 dig_ctrl_inst.latch_mem_inst.RAM\[62\]\[0\]
+ sky130_fd_sc_hd__and3_2
X_2203_ VGND VDPWR VDPWR VGND _0890_ _0892_ _0891_ sky130_fd_sc_hd__and2b_1
X_2134_ VDPWR VGND VDPWR VGND _0825_ dig_ctrl_inst.cpu_inst.data\[1\] _0743_ _0826_
+ net164 sky130_fd_sc_hd__a22o_1
X_2065_ VGND VDPWR VDPWR VGND _0758_ net300 _0755_ _0757_ _0199_ sky130_fd_sc_hd__o211a_1
X_1849_ VDPWR VGND VDPWR VGND _0131_ dig_ctrl_inst.latch_mem_inst.RAM\[1\]\[4\] _1130_
+ _0557_ dig_ctrl_inst.latch_mem_inst.RAM\[29\]\[4\] sky130_fd_sc_hd__a22o_1
X_1918_ VDPWR VGND VDPWR VGND _0624_ net68 net111 dig_ctrl_inst.latch_mem_inst.RAM\[18\]\[6\]
+ sky130_fd_sc_hd__and3_2
XFILLER_0_39_137 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_54_118 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[55\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[55\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[55\] clknet_leaf_17_clk sky130_fd_sc_hd__dlclkp_1
X_1703_ VDPWR VGND VDPWR VGND _0413_ net73 net123 dig_ctrl_inst.latch_mem_inst.RAM\[14\]\[2\]
+ sky130_fd_sc_hd__and3_2
Xclkbuf_leaf_11_clk VGND VDPWR VDPWR VGND clknet_leaf_11_clk clknet_1_0__leaf_clk
+ sky130_fd_sc_hd__clkbuf_8
X_1634_ VGND VDPWR VDPWR VGND _0345_ net43 net80 net115 dig_ctrl_inst.latch_mem_inst.RAM\[61\]\[1\]
+ sky130_fd_sc_hd__and4_1
X_1565_ VDPWR VGND VDPWR VGND net125 net97 _0277_ sky130_fd_sc_hd__and2_2
X_1496_ VGND VDPWR VDPWR VGND _0213_ dig_ctrl_inst.cpu_inst.data\[2\] _0198_ _1060_
+ sky130_fd_sc_hd__mux2_1
X_2048_ VGND VDPWR VDPWR VGND _0044_ net354 _0161_ dig_ctrl_inst.cpu_inst.cpu_state\[2\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_3 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2117_ VGND VDPWR VDPWR VGND net157 _0760_ _0258_ _0766_ _0809_ sky130_fd_sc_hd__o22a_1
Xfanout69 VDPWR VGND VDPWR VGND net69 net71 sky130_fd_sc_hd__buf_2
Xfanout58 VDPWR VGND VDPWR VGND net58 net59 sky130_fd_sc_hd__buf_2
XFILLER_0_17_310 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
Xfanout47 VGND VDPWR VDPWR VGND _0147_ net47 sky130_fd_sc_hd__clkbuf_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[62\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[62\]\[6\] net195 dig_ctrl_inst.latch_mem_inst.gclk\[62\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[58\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[58\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[58\] sky130_fd_sc_hd__clkbuf_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[51\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[51\]\[4\] net212 dig_ctrl_inst.latch_mem_inst.gclk\[51\]
+ sky130_fd_sc_hd__dlxtp_1
Xclkload17 VGND VDPWR VDPWR VGND clkload17/Y clknet_leaf_19_clk sky130_fd_sc_hd__inv_12
X_1350_ VGND VDPWR VDPWR VGND _0132_ net106 net82 net69 sky130_fd_sc_hd__and3_4
X_1281_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[0\] net121 net152
+ net130 sky130_fd_sc_hd__and3_2
Xclkbuf_leaf_0_clk VGND VDPWR VDPWR VGND clknet_leaf_0_clk clknet_1_1__leaf_clk sky130_fd_sc_hd__clkbuf_8
Xdig_ctrl_inst.latch_mem_inst.gen_words\[40\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[40\]\[2\] net224 dig_ctrl_inst.latch_mem_inst.gclk\[40\]
+ sky130_fd_sc_hd__dlxtp_1
Xfanout204 VGND VDPWR VDPWR VGND net206 net204 sky130_fd_sc_hd__clkbuf_2
X_1617_ VDPWR VGND VDPWR VGND _0148_ dig_ctrl_inst.latch_mem_inst.RAM\[44\]\[0\] _0144_
+ _0329_ dig_ctrl_inst.latch_mem_inst.RAM\[49\]\[0\] sky130_fd_sc_hd__a22o_1
XFILLER_0_41_132 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_1_295 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
Xfanout248 VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.cpu_state\[0\] net248 sky130_fd_sc_hd__clkbuf_4
Xfanout237 VGND VDPWR VDPWR VGND net238 net237 sky130_fd_sc_hd__clkbuf_2
Xfanout226 VGND VDPWR VDPWR VGND net227 net226 sky130_fd_sc_hd__clkbuf_2
X_1548_ VDPWR VGND VDPWR VGND _0261_ _0258_ _0260_ sky130_fd_sc_hd__and2_1
Xfanout215 VGND VDPWR VDPWR VGND net216 net215 sky130_fd_sc_hd__clkbuf_2
X_1479_ VDPWR VGND VDPWR VGND _0198_ net285 _1031_ sky130_fd_sc_hd__or2_2
Xfanout259 VDPWR VGND VDPWR VGND net259 dig_ctrl_inst.cpu_inst.arg1\[0\] sky130_fd_sc_hd__buf_2
XFILLER_0_20_338 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_1_3 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_29 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[55\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[55\]\[5\] net203 dig_ctrl_inst.latch_mem_inst.gclk\[55\]
+ sky130_fd_sc_hd__dlxtp_1
X_1402_ VDPWR VGND VDPWR VGND _0156_ net49 net92 net107 sky130_fd_sc_hd__and3_2
X_2520_ VDPWR VGND VDPWR VGND uio_oe[1] net270 sky130_fd_sc_hd__buf_2
XFILLER_0_23_165 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2451_ VGND VDPWR VDPWR VGND clknet_leaf_10_clk _0059_ net142 dig_ctrl_inst.cpu_inst.r1\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_2382_ VGND VDPWR VDPWR VGND clknet_leaf_3_clk net8 net175 dig_ctrl_inst.synchronizer_port_i_inst\[5\].pipe\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_1264_ VGND VDPWR VDPWR VGND _1105_ _1111_ _1002_ _1112_ _1098_ dig_ctrl_inst.spi_addr\[5\]
+ sky130_fd_sc_hd__o32a_4
Xinput4 VGND VDPWR VDPWR VGND net4 ui_in[1] sky130_fd_sc_hd__clkbuf_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[44\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[44\]\[3\] net221 dig_ctrl_inst.latch_mem_inst.gclk\[44\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_36_41 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
X_1333_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[21\] net150 _0124_
+ sky130_fd_sc_hd__and2_1
X_1195_ VGND VDPWR VDPWR VGND net264 _1043_ dig_ctrl_inst.cpu_inst.r1\[3\] sky130_fd_sc_hd__and2b_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[33\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[33\]\[1\] net233 dig_ctrl_inst.latch_mem_inst.gclk\[33\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[10\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[10\]\[6\] net195 dig_ctrl_inst.latch_mem_inst.gclk\[10\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[59\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[59\]\[6\] net195 dig_ctrl_inst.latch_mem_inst.gclk\[59\]
+ sky130_fd_sc_hd__dlxtp_1
X_1951_ VDPWR VGND VDPWR VGND _0657_ net43 net96 dig_ctrl_inst.latch_mem_inst.RAM\[52\]\[6\]
+ sky130_fd_sc_hd__and3_2
X_1882_ VGND VDPWR VDPWR VGND _0589_ net63 net100 net103 dig_ctrl_inst.latch_mem_inst.RAM\[23\]\[5\]
+ sky130_fd_sc_hd__and4_1
X_2503_ VGND VDPWR VDPWR VGND clknet_leaf_5_clk _0100_ net177 net33 sky130_fd_sc_hd__dfrtp_1
X_2434_ VDPWR VGND VDPWR VGND clknet_leaf_8_clk net347 dig_ctrl_inst.cpu_inst.prev_state\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[48\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[48\]\[4\] net323 dig_ctrl_inst.latch_mem_inst.gclk\[48\]
+ sky130_fd_sc_hd__dlxtp_1
X_2365_ VDPWR VGND VDPWR VGND _0992_ _0623_ _0565_ _0506_ sky130_fd_sc_hd__and3_2
XFILLER_0_11_113 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1316_ VDPWR VGND VDPWR VGND _0115_ _1047_ net135 _1093_ _1077_ _1075_ sky130_fd_sc_hd__o2111a_1
X_1247_ VDPWR VGND VDPWR VGND _1047_ net135 _1093_ _1076_ _1095_ _1078_ sky130_fd_sc_hd__a2111oi_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[37\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[37\]\[2\] net228 dig_ctrl_inst.latch_mem_inst.gclk\[37\]
+ sky130_fd_sc_hd__dlxtp_1
X_1178_ VGND VDPWR VDPWR VGND _1011_ _1026_ _1015_ net283 _1019_ net298 sky130_fd_sc_hd__o32ai_4
X_2296_ VGND VDPWR VDPWR VGND _0059_ _0974_ _0967_ net361 sky130_fd_sc_hd__mux2_1
XANTENNA_31 VGND VDPWR VDPWR VGND net19 sky130_fd_sc_hd__diode_2
XANTENNA_20 VGND VDPWR VDPWR VGND net100 sky130_fd_sc_hd__diode_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[26\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[26\]\[0\] net246 dig_ctrl_inst.latch_mem_inst.gclk\[26\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_69_113 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
Xdig_ctrl_inst.latch_mem_inst.gen_words\[14\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[14\]\[7\] net185 dig_ctrl_inst.latch_mem_inst.gclk\[14\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_0_305 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2081_ VGND VDPWR VDPWR VGND _0763_ _0765_ _0773_ _0774_ sky130_fd_sc_hd__o21a_1
X_2150_ VDPWR VGND VDPWR VGND _0838_ _0839_ _0841_ _0840_ net167 net170 sky130_fd_sc_hd__a221o_1
X_1934_ VGND VDPWR VDPWR VGND _0640_ net68 net118 net132 dig_ctrl_inst.latch_mem_inst.RAM\[17\]\[6\]
+ sky130_fd_sc_hd__and4_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[8\].gen_latches\[0\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[8\]\[0\] net242 dig_ctrl_inst.latch_mem_inst.gclk\[8\]
+ sky130_fd_sc_hd__dlxtp_1
X_1796_ VDPWR VGND VDPWR VGND _0505_ net39 _0504_ _0288_ dig_ctrl_inst.latch_mem_inst.RAM\[0\]\[3\]
+ sky130_fd_sc_hd__o2bb2a_1
X_1865_ VDPWR VGND VDPWR VGND _0572_ net83 net124 dig_ctrl_inst.latch_mem_inst.RAM\[10\]\[5\]
+ sky130_fd_sc_hd__and3_2
X_2348_ VGND VDPWR VDPWR VGND _0098_ net31 _0987_ dig_ctrl_inst.cpu_inst.port_o\[3\]
+ sky130_fd_sc_hd__mux2_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[62\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[62\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[62\] clknet_leaf_0_clk sky130_fd_sc_hd__dlclkp_1
X_2417_ VGND VDPWR VDPWR VGND clknet_leaf_10_clk _0025_ net140 dig_ctrl_inst.cpu_inst.skip
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_10_Left_88 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2279_ VDPWR VGND VDPWR VGND dig_ctrl_inst.spi_data_o\[7\] _0804_ _0965_ dig_ctrl_inst.synchronizer_port_i_inst\[7\].out
+ _0802_ sky130_fd_sc_hd__a22oi_2
Xhold109 VGND VDPWR VDPWR VGND net391 dig_ctrl_inst.spi_receiver_inst.spi_cnt\[2\]
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_333 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1581_ VGND VDPWR VDPWR VGND _0293_ net48 net82 net118 dig_ctrl_inst.latch_mem_inst.RAM\[61\]\[0\]
+ sky130_fd_sc_hd__and4_1
X_1650_ VDPWR VGND VDPWR VGND _0361_ net42 net109 dig_ctrl_inst.latch_mem_inst.RAM\[50\]\[1\]
+ sky130_fd_sc_hd__and3_2
X_2202_ VGND VDPWR VDPWR VGND net159 _0891_ _0867_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_146 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_0_113 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_44_41 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2133_ VGND VDPWR VDPWR VGND _1019_ _0825_ _1015_ sky130_fd_sc_hd__nor2_2
X_2064_ VDPWR VGND VDPWR VGND _1024_ _1020_ _0756_ _0757_ sky130_fd_sc_hd__a21o_1
X_1917_ VGND VDPWR VDPWR VGND _0031_ _0622_ _0276_ net252 sky130_fd_sc_hd__mux2_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[8\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[8\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[8\] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_71 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1848_ VDPWR VGND VDPWR VGND _0155_ dig_ctrl_inst.latch_mem_inst.RAM\[9\]\[4\] _1143_
+ _0556_ dig_ctrl_inst.latch_mem_inst.RAM\[58\]\[4\] sky130_fd_sc_hd__a22o_1
X_1779_ VDPWR VGND VDPWR VGND _0488_ net56 net72 dig_ctrl_inst.latch_mem_inst.RAM\[46\]\[3\]
+ sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[22\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[22\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[22\] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_62_141 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1564_ VDPWR VGND VDPWR VGND net182 _0200_ _0276_ sky130_fd_sc_hd__and2_2
X_1633_ VGND VDPWR VDPWR VGND _0344_ net42 net90 net102 dig_ctrl_inst.latch_mem_inst.RAM\[59\]\[1\]
+ sky130_fd_sc_hd__and4_1
X_1702_ VDPWR VGND VDPWR VGND _0412_ net46 net130 dig_ctrl_inst.latch_mem_inst.RAM\[48\]\[2\]
+ sky130_fd_sc_hd__and3_2
X_1495_ VDPWR VGND VDPWR VGND _0212_ _0210_ dig_ctrl_inst.cpu_inst.ip\[1\] dig_ctrl_inst.cpu_inst.ip\[0\]
+ sky130_fd_sc_hd__and3_2
X_2047_ VGND VDPWR VDPWR VGND _0043_ net349 _0161_ dig_ctrl_inst.cpu_inst.cpu_state\[1\]
+ sky130_fd_sc_hd__mux2_1
X_2116_ VGND VDPWR VDPWR VGND _0808_ _0776_ net157 _0761_ sky130_fd_sc_hd__mux2_1
Xfanout59 VDPWR VGND VDPWR VGND net60 net59 sky130_fd_sc_hd__buf_4
Xfanout48 VDPWR VGND VDPWR VGND net49 net48 sky130_fd_sc_hd__buf_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[63\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[63\]\[1\] net237 dig_ctrl_inst.latch_mem_inst.gclk\[63\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_44_141 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_17_322 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_13_Left_91 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_27_108 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1280_ VGND VDPWR VDPWR VGND _1112_ _1127_ _1128_ sky130_fd_sc_hd__nor2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[40\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[40\]\[6\] net196 dig_ctrl_inst.latch_mem_inst.gclk\[40\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_25_10 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
Xfanout238 VGND VDPWR VDPWR VGND net239 net238 sky130_fd_sc_hd__clkbuf_2
Xfanout205 VGND VDPWR VDPWR VGND net205 net206 sky130_fd_sc_hd__buf_1
X_1616_ VGND VDPWR VDPWR VGND _0122_ dig_ctrl_inst.latch_mem_inst.RAM\[19\]\[0\] _0293_
+ _0294_ _0302_ _0328_ sky130_fd_sc_hd__a2111o_1
Xfanout216 VDPWR VGND VDPWR VGND net216 net329 sky130_fd_sc_hd__buf_2
X_1547_ VGND VDPWR VDPWR VGND _0260_ net158 net164 sky130_fd_sc_hd__or2_1
Xfanout227 VGND VDPWR VDPWR VGND net231 net227 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_5_31 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
Xfanout249 VGND VDPWR VDPWR VGND net251 net249 sky130_fd_sc_hd__clkbuf_4
X_1478_ VGND VDPWR VDPWR VGND _0018_ dig_ctrl_inst.cpu_inst.port_o\[7\] _0176_ dig_ctrl_inst.cpu_inst.r0\[7\]
+ sky130_fd_sc_hd__mux2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[56\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[56\]\[0\] net242 dig_ctrl_inst.latch_mem_inst.gclk\[56\]
+ sky130_fd_sc_hd__dlxtp_1
X_2381_ VGND VDPWR VDPWR VGND clknet_leaf_4_clk net338 net174 dig_ctrl_inst.synchronizer_port_i_inst\[6\].out
+ sky130_fd_sc_hd__dfrtp_1
X_2450_ VGND VDPWR VDPWR VGND clknet_leaf_7_clk _0058_ net144 dig_ctrl_inst.cpu_inst.r1\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_1401_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[58\] net50 net85
+ net155 sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[0\].gen_latches\[2\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[0\]\[2\] net226 dig_ctrl_inst.latch_mem_inst.gclk\[0\]
+ sky130_fd_sc_hd__dlxtp_1
Xinput5 VGND VDPWR VDPWR VGND net5 ui_in[2] sky130_fd_sc_hd__clkbuf_1
X_1194_ VGND VDPWR VDPWR VGND net267 _1042_ dig_ctrl_inst.cpu_inst.r2\[3\] sky130_fd_sc_hd__and2b_1
X_1263_ VDPWR VGND VDPWR VGND _1110_ _1039_ net249 _1111_ sky130_fd_sc_hd__a21o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[44\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[44\]\[7\] net189 dig_ctrl_inst.latch_mem_inst.gclk\[44\]
+ sky130_fd_sc_hd__dlxtp_1
X_1332_ VDPWR VGND VDPWR VGND _0124_ net62 net99 net116 sky130_fd_sc_hd__and3_2
XFILLER_0_52_85 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[15\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[15\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[15\] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_72_3 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[33\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[33\]\[5\] net201 dig_ctrl_inst.latch_mem_inst.gclk\[33\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[22\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[22\]\[3\] net220 dig_ctrl_inst.latch_mem_inst.gclk\[22\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[11\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[11\]\[1\] net238 dig_ctrl_inst.latch_mem_inst.gclk\[11\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_29_Left_107 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_38_Left_116 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1950_ VDPWR VGND VDPWR VGND _0656_ net57 net88 dig_ctrl_inst.latch_mem_inst.RAM\[40\]\[6\]
+ sky130_fd_sc_hd__and3_2
XFILLER_0_22_22 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
X_2502_ VGND VDPWR VDPWR VGND clknet_leaf_5_clk _0099_ net177 net32 sky130_fd_sc_hd__dfrtp_1
X_1881_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[1\]\[5\] _1130_ _0588_
+ _0152_ dig_ctrl_inst.latch_mem_inst.RAM\[54\]\[5\] _0587_ sky130_fd_sc_hd__a221o_1
XFILLER_0_22_99 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_3_325 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_2364_ VGND VDPWR VDPWR VGND _0338_ _0991_ _0623_ _0506_ _0398_ sky130_fd_sc_hd__o211ai_1
X_1315_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[13\] net155 _0114_
+ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_47_Left_125 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[4\].gen_latches\[3\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[4\]\[3\] net220 dig_ctrl_inst.latch_mem_inst.gclk\[4\]
+ sky130_fd_sc_hd__dlxtp_1
X_2433_ VGND VDPWR VDPWR VGND clknet_leaf_13_clk _0041_ net139 dig_ctrl_inst.cpu_inst.data\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_1246_ VGND VDPWR VDPWR VGND net249 _1079_ _1091_ _1085_ _1094_ _1092_ sky130_fd_sc_hd__o41ai_2
XPHY_EDGE_ROW_56_Left_134 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1177_ VGND VDPWR VDPWR VGND _1019_ _1017_ _1011_ _1025_ net181 _1015_ sky130_fd_sc_hd__o32a_4
X_2295_ VGND VDPWR VDPWR VGND _0946_ _0943_ _0974_ _0751_ sky130_fd_sc_hd__o21ai_1
XANTENNA_21 VGND VDPWR VDPWR VGND net329 sky130_fd_sc_hd__diode_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[37\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[37\]\[6\] net195 dig_ctrl_inst.latch_mem_inst.gclk\[37\]
+ sky130_fd_sc_hd__dlxtp_1
XANTENNA_32 VGND VDPWR VDPWR VGND _1135_ sky130_fd_sc_hd__diode_2
XANTENNA_10 VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[19\] sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_65_Left_143 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_74_Left_152 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[26\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[26\]\[4\] net211 dig_ctrl_inst.latch_mem_inst.gclk\[26\]
+ sky130_fd_sc_hd__dlxtp_1
Xmax_cap89 VGND VDPWR VDPWR VGND net89 _1141_ sky130_fd_sc_hd__buf_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[15\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[15\]\[2\] net229 dig_ctrl_inst.latch_mem_inst.gclk\[15\]
+ sky130_fd_sc_hd__dlxtp_1
X_2080_ VGND VDPWR VDPWR VGND _0773_ _0767_ _0768_ _0771_ _0772_ sky130_fd_sc_hd__o211a_1
X_1933_ VDPWR VGND VDPWR VGND _0639_ net76 net122 dig_ctrl_inst.latch_mem_inst.RAM\[12\]\[6\]
+ sky130_fd_sc_hd__and3_2
X_1864_ VDPWR VGND VDPWR VGND _0571_ net49 net88 dig_ctrl_inst.latch_mem_inst.RAM\[56\]\[5\]
+ sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[8\].gen_latches\[4\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[8\]\[4\] net209 dig_ctrl_inst.latch_mem_inst.gclk\[8\]
+ sky130_fd_sc_hd__dlxtp_1
X_1795_ VGND VDPWR VDPWR VGND _0504_ _0503_ _0486_ _0469_ _0464_ sky130_fd_sc_hd__nor4_1
X_2347_ VGND VDPWR VDPWR VGND _0097_ net30 _0987_ dig_ctrl_inst.cpu_inst.port_o\[2\]
+ sky130_fd_sc_hd__mux2_1
X_2416_ VGND VDPWR VDPWR VGND clknet_leaf_13_clk _0024_ net140 dig_ctrl_inst.cpu_inst.ip\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_2278_ VDPWR VGND VDPWR VGND _0233_ _0964_ _0944_ sky130_fd_sc_hd__xor2_1
X_1229_ VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_addr\[0\] _1002_ _1077_ sky130_fd_sc_hd__nor2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[19\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[19\]\[3\] net215 dig_ctrl_inst.latch_mem_inst.gclk\[19\]
+ sky130_fd_sc_hd__dlxtp_1
X_1580_ VDPWR VGND VDPWR VGND _0292_ net66 net87 dig_ctrl_inst.latch_mem_inst.RAM\[24\]\[0\]
+ sky130_fd_sc_hd__and3_2
XFILLER_0_0_103 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_0_169 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_2132_ VGND VDPWR VDPWR VGND _0793_ _0254_ _0785_ _0255_ _0824_ _0823_ sky130_fd_sc_hd__o221a_1
X_2201_ VGND VDPWR VDPWR VGND net159 _0867_ _0890_ sky130_fd_sc_hd__nor2_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[61\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[61\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[61\] sky130_fd_sc_hd__clkbuf_4
X_2063_ VGND VDPWR VDPWR VGND _0753_ _0751_ _0756_ sky130_fd_sc_hd__or2_4
XFILLER_0_63_109 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1847_ VGND VDPWR VDPWR VGND _0156_ dig_ctrl_inst.latch_mem_inst.RAM\[59\]\[4\] _0552_
+ _0553_ _0554_ _0555_ sky130_fd_sc_hd__a2111o_1
X_1916_ VGND VDPWR VDPWR VGND net37 net36 _0288_ dig_ctrl_inst.latch_mem_inst.RAM\[0\]\[5\]
+ _0623_ sky130_fd_sc_hd__a2bb2o_1
X_1778_ VDPWR VGND VDPWR VGND _0487_ net56 net129 dig_ctrl_inst.latch_mem_inst.RAM\[32\]\[3\]
+ sky130_fd_sc_hd__and3_2
XFILLER_0_35_312 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1701_ VDPWR VGND VDPWR VGND _0411_ net50 net111 dig_ctrl_inst.latch_mem_inst.RAM\[50\]\[2\]
+ sky130_fd_sc_hd__and3_2
XFILLER_0_39_20 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_337 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2523__272 VGND VDPWR VDPWR VGND net272 _2523__272/HI sky130_fd_sc_hd__conb_1
X_1632_ VDPWR VGND VDPWR VGND _0343_ net67 net94 dig_ctrl_inst.latch_mem_inst.RAM\[22\]\[1\]
+ sky130_fd_sc_hd__and3_2
X_1563_ VDPWR VGND VDPWR VGND _0274_ dig_ctrl_inst.cpu_inst.skip _0174_ _0025_ _0275_
+ sky130_fd_sc_hd__a22o_1
X_1494_ VGND VDPWR VDPWR VGND _0211_ _0204_ _0210_ sky130_fd_sc_hd__or2_1
X_2115_ VGND VDPWR VDPWR VGND _0045_ _0807_ net41 dig_ctrl_inst.cpu_inst.r0\[0\] sky130_fd_sc_hd__mux2_1
Xfanout49 VDPWR VGND VDPWR VGND net50 net49 sky130_fd_sc_hd__buf_4
X_2046_ VGND VDPWR VDPWR VGND _0042_ net346 _0161_ dig_ctrl_inst.cpu_inst.cpu_state\[0\]
+ sky130_fd_sc_hd__mux2_1
X_2530__276 VGND VDPWR VDPWR VGND net276 _2530__276/HI sky130_fd_sc_hd__conb_1
XFILLER_0_36_109 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_44_197 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[63\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[63\]\[5\] net203 dig_ctrl_inst.latch_mem_inst.gclk\[63\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[52\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[52\]\[3\] net216 dig_ctrl_inst.latch_mem_inst.gclk\[52\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_35_120 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[41\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[41\]\[1\] net236 dig_ctrl_inst.latch_mem_inst.gclk\[41\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_23_337 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_26_153 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_26_197 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1477_ VGND VDPWR VDPWR VGND _0017_ dig_ctrl_inst.cpu_inst.port_o\[6\] _0176_ dig_ctrl_inst.cpu_inst.r0\[6\]
+ sky130_fd_sc_hd__mux2_1
Xfanout239 VGND VDPWR VDPWR VGND net327 net239 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_41_189 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xfanout206 VGND VDPWR VDPWR VGND net206 net207 sky130_fd_sc_hd__buf_1
Xfanout228 VGND VDPWR VDPWR VGND net231 net228 sky130_fd_sc_hd__clkbuf_2
X_1615_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[12\]\[0\] _1148_ _0327_
+ _0278_ dig_ctrl_inst.latch_mem_inst.RAM\[5\]\[0\] _0289_ sky130_fd_sc_hd__a221o_1
XFILLER_0_1_275 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xfanout217 VGND VDPWR VDPWR VGND net219 net217 sky130_fd_sc_hd__clkbuf_2
X_1546_ VGND VDPWR VDPWR VGND net158 net164 _0259_ sky130_fd_sc_hd__nor2_1
X_2029_ VDPWR VGND VDPWR VGND _0733_ _0732_ _0731_ _0730_ _0734_ sky130_fd_sc_hd__or4_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[56\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[56\]\[4\] net214 dig_ctrl_inst.latch_mem_inst.gclk\[56\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_11_57 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[45\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[45\]\[2\] net224 dig_ctrl_inst.latch_mem_inst.gclk\[45\]
+ sky130_fd_sc_hd__dlxtp_1
X_2380_ VGND VDPWR VDPWR VGND clknet_leaf_3_clk net9 net175 dig_ctrl_inst.synchronizer_port_i_inst\[6\].pipe\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_1400_ VDPWR VGND VDPWR VGND net83 _0147_ _0155_ sky130_fd_sc_hd__and2_2
X_1331_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[20\] net68 net97
+ net156 sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[54\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[54\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[54\] sky130_fd_sc_hd__clkbuf_4
Xinput6 VGND VDPWR VDPWR VGND net6 ui_in[3] sky130_fd_sc_hd__clkbuf_1
X_1193_ VDPWR VGND VDPWR VGND _1041_ dig_ctrl_inst.cpu_inst.r3\[3\] net264 net267
+ sky130_fd_sc_hd__and3_2
X_1262_ VGND VDPWR VDPWR VGND net181 _1106_ _1107_ _1108_ _1109_ _1110_ sky130_fd_sc_hd__o41a_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[34\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[34\]\[0\] net245 dig_ctrl_inst.latch_mem_inst.gclk\[34\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[0\].gen_latches\[6\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[0\]\[6\] net193 dig_ctrl_inst.latch_mem_inst.gclk\[0\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_6_323 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_1529_ VGND VDPWR VDPWR VGND _1103_ _0242_ net160 sky130_fd_sc_hd__nand2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[22\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[22\]\[7\] net184 dig_ctrl_inst.latch_mem_inst.gclk\[22\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_14_Right_14 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[11\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[11\]\[5\] net204 dig_ctrl_inst.latch_mem_inst.gclk\[11\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_23_Right_23 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1880_ VDPWR VGND VDPWR VGND _0587_ net60 net86 dig_ctrl_inst.latch_mem_inst.RAM\[40\]\[5\]
+ sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[49\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[49\]\[3\] net217 dig_ctrl_inst.latch_mem_inst.gclk\[49\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_32_Right_32 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2501_ VGND VDPWR VDPWR VGND clknet_leaf_5_clk _0098_ net178 net31 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_337 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1314_ VGND VDPWR VDPWR VGND _0114_ net126 net119 net82 sky130_fd_sc_hd__and3_4
X_2363_ VGND VDPWR VDPWR VGND _0201_ _0990_ _0989_ sky130_fd_sc_hd__nand2_1
X_2294_ VGND VDPWR VDPWR VGND _0058_ _0973_ _0967_ net365 sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_41_Right_41 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[4\].gen_latches\[7\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[4\]\[7\] net187 dig_ctrl_inst.latch_mem_inst.gclk\[4\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[38\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[38\]\[1\] net234 dig_ctrl_inst.latch_mem_inst.gclk\[38\]
+ sky130_fd_sc_hd__dlxtp_1
X_2432_ VGND VDPWR VDPWR VGND clknet_leaf_13_clk _0040_ net139 dig_ctrl_inst.cpu_inst.data\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_1245_ VGND VDPWR VDPWR VGND _1093_ _1092_ _1085_ _1091_ net289 net249 sky130_fd_sc_hd__o41a_4
XPHY_EDGE_ROW_50_Right_50 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1176_ VDPWR VGND VDPWR VGND _1024_ _0998_ net264 sky130_fd_sc_hd__and2_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[13\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[13\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[13\] clknet_leaf_2_clk sky130_fd_sc_hd__dlclkp_1
XANTENNA_33 VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.port_o\[5\] sky130_fd_sc_hd__diode_2
XANTENNA_22 VGND VDPWR VDPWR VGND net322 sky130_fd_sc_hd__diode_2
XANTENNA_11 VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[32\] sky130_fd_sc_hd__diode_2
XFILLER_0_10_192 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[15\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[15\]\[6\] net191 dig_ctrl_inst.latch_mem_inst.gclk\[15\]
+ sky130_fd_sc_hd__dlxtp_1
X_1863_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[27\]\[5\] _0130_ _0570_
+ _0278_ dig_ctrl_inst.latch_mem_inst.RAM\[5\]\[5\] _0569_ sky130_fd_sc_hd__a221o_1
X_1932_ VDPWR VGND VDPWR VGND _0638_ net83 net124 dig_ctrl_inst.latch_mem_inst.RAM\[10\]\[6\]
+ sky130_fd_sc_hd__and3_2
X_2526__281 VGND VDPWR VDPWR VGND _2526__281/LO net281 sky130_fd_sc_hd__conb_1
X_2415_ VGND VDPWR VDPWR VGND clknet_leaf_13_clk _0023_ net140 dig_ctrl_inst.cpu_inst.ip\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_1794_ VDPWR VGND VDPWR VGND _0494_ _0502_ _0498_ _0490_ _0503_ sky130_fd_sc_hd__or4_1
X_2346_ VGND VDPWR VDPWR VGND _0096_ net389 _0987_ dig_ctrl_inst.cpu_inst.port_o\[1\]
+ sky130_fd_sc_hd__mux2_1
X_1228_ VDPWR VGND VDPWR VGND _1074_ _1030_ _1067_ dig_ctrl_inst.cpu_inst.ip\[0\]
+ _1028_ _1076_ sky130_fd_sc_hd__a221o_2
XFILLER_0_58_85 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_28_3 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2277_ VGND VDPWR VDPWR VGND _0788_ _0951_ _0962_ _0963_ sky130_fd_sc_hd__o21a_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[19\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[19\]\[7\] net188 dig_ctrl_inst.latch_mem_inst.gclk\[19\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[47\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[47\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[47\] sky130_fd_sc_hd__clkbuf_4
X_2062_ VGND VDPWR VDPWR VGND _0751_ _0753_ _0755_ sky130_fd_sc_hd__nor2_1
X_2131_ VGND VDPWR VDPWR VGND _0823_ _0791_ net163 _0786_ sky130_fd_sc_hd__mux2_1
X_2200_ VDPWR VGND VDPWR VGND net167 _0771_ _0889_ _0781_ _0888_ net170 sky130_fd_sc_hd__a221o_1
XFILLER_0_44_98 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_60_97 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_1846_ VDPWR VGND VDPWR VGND _0554_ net49 net88 dig_ctrl_inst.latch_mem_inst.RAM\[56\]\[4\]
+ sky130_fd_sc_hd__and3_2
X_1777_ VDPWR VGND VDPWR VGND _0477_ _0485_ _0481_ _0473_ _0486_ sky130_fd_sc_hd__or4_1
X_1915_ VDPWR VGND VDPWR VGND _0622_ net37 net36 _0288_ dig_ctrl_inst.latch_mem_inst.RAM\[0\]\[5\]
+ sky130_fd_sc_hd__o2bb2a_1
XPHY_EDGE_ROW_4_Right_4 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2329_ VGND VDPWR VDPWR VGND _0081_ dig_ctrl_inst.spi_data_o\[2\] _0180_ dig_ctrl_inst.spi_data_o\[1\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_132 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
Xclone12 VGND VDPWR VDPWR VGND net294 _1144_ sky130_fd_sc_hd__clkbuf_1
X_1700_ VDPWR VGND VDPWR VGND _0410_ net49 net85 dig_ctrl_inst.latch_mem_inst.RAM\[58\]\[2\]
+ sky130_fd_sc_hd__and3_2
X_1631_ VDPWR VGND VDPWR VGND _0342_ net67 net76 dig_ctrl_inst.latch_mem_inst.RAM\[28\]\[1\]
+ sky130_fd_sc_hd__and3_2
XFILLER_0_30_34 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_30_23 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_39_32 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_3_clk VGND VDPWR VDPWR VGND clknet_leaf_3_clk clknet_1_1__leaf_clk sky130_fd_sc_hd__clkbuf_8
X_1493_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.ip\[2\] dig_ctrl_inst.cpu_inst.ip\[1\]
+ dig_ctrl_inst.cpu_inst.ip\[0\] _0210_ _0173_ sky130_fd_sc_hd__a31oi_1
X_1562_ VDPWR VGND VDPWR VGND _0275_ _0175_ dig_ctrl_inst.cpu_inst.instr\[7\] dig_ctrl_inst.cpu_inst.instr\[6\]
+ sky130_fd_sc_hd__and3_2
X_2114_ VGND VDPWR VDPWR VGND _0798_ _0807_ _0806_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_53 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2045_ VGND VDPWR VDPWR VGND _0041_ _0740_ _0741_ net387 sky130_fd_sc_hd__mux2_1
X_1829_ VGND VDPWR VDPWR VGND _0537_ net51 net90 net114 dig_ctrl_inst.latch_mem_inst.RAM\[41\]\[4\]
+ sky130_fd_sc_hd__and4_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[4\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[4\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[4\] sky130_fd_sc_hd__clkbuf_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[52\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[52\]\[7\] net190 dig_ctrl_inst.latch_mem_inst.gclk\[52\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[41\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[41\]\[5\] net199 dig_ctrl_inst.latch_mem_inst.gclk\[41\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[30\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[30\]\[3\] net222 dig_ctrl_inst.latch_mem_inst.gclk\[30\]
+ sky130_fd_sc_hd__dlxtp_1
X_1614_ VDPWR VGND VDPWR VGND _0318_ _0325_ _0313_ _0326_ sky130_fd_sc_hd__or3_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[18\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[18\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[18\] clknet_leaf_17_clk sky130_fd_sc_hd__dlclkp_1
Xfanout218 VGND VDPWR VDPWR VGND net218 net219 sky130_fd_sc_hd__buf_1
Xfanout229 VGND VDPWR VDPWR VGND net230 net229 sky130_fd_sc_hd__clkbuf_2
X_1476_ VGND VDPWR VDPWR VGND _0016_ dig_ctrl_inst.cpu_inst.port_o\[5\] _0176_ dig_ctrl_inst.cpu_inst.r0\[5\]
+ sky130_fd_sc_hd__mux2_1
Xfanout207 VGND VDPWR VDPWR VGND net326 net207 sky130_fd_sc_hd__clkbuf_2
X_1545_ VGND VDPWR VDPWR VGND _1066_ _0258_ _1019_ dig_ctrl_inst.cpu_inst.r0\[0\]
+ _1065_ net165 sky130_fd_sc_hd__o221ai_4
XFILLER_0_1_254 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_5_99 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2028_ VDPWR VGND VDPWR VGND _0149_ dig_ctrl_inst.latch_mem_inst.RAM\[13\]\[7\] _0114_
+ _0733_ dig_ctrl_inst.latch_mem_inst.RAM\[51\]\[7\] sky130_fd_sc_hd__a22o_1
XFILLER_0_10_3 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_17_165 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[20\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[20\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[20\] clknet_leaf_19_clk sky130_fd_sc_hd__dlclkp_1
X_1261_ VDPWR VGND VDPWR VGND net263 dig_ctrl_inst.cpu_inst.r0\[5\] net267 _1109_
+ sky130_fd_sc_hd__or3_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[45\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[45\]\[6\] net197 dig_ctrl_inst.latch_mem_inst.gclk\[45\]
+ sky130_fd_sc_hd__dlxtp_1
X_1330_ VDPWR VGND VDPWR VGND _0123_ net97 net68 sky130_fd_sc_hd__and2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[1\].gen_latches\[1\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[1\]\[1\] net237 dig_ctrl_inst.latch_mem_inst.gclk\[1\]
+ sky130_fd_sc_hd__dlxtp_1
Xinput7 VGND VDPWR VDPWR VGND net7 ui_in[4] sky130_fd_sc_hd__clkbuf_1
X_1192_ VDPWR VGND VDPWR VGND dig_ctrl_inst.cpu_inst.cpu_state\[1\] _0999_ net248
+ _1040_ sky130_fd_sc_hd__or3_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[34\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[34\]\[4\] net213 dig_ctrl_inst.latch_mem_inst.gclk\[34\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_6_335 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
Xdig_ctrl_inst.latch_mem_inst.gen_words\[23\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[23\]\[2\] net225 dig_ctrl_inst.latch_mem_inst.gclk\[23\]
+ sky130_fd_sc_hd__dlxtp_1
X_1459_ VGND VDPWR VDPWR VGND _0190_ _0185_ dig_ctrl_inst.spi_addr\[1\] dig_ctrl_inst.spi_addr\[0\]
+ dig_ctrl_inst.spi_addr\[2\] sky130_fd_sc_hd__a31o_1
X_1528_ VDPWR VGND VDPWR VGND _0241_ _1103_ net160 sky130_fd_sc_hd__and2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[12\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[12\]\[0\] net243 dig_ctrl_inst.latch_mem_inst.gclk\[12\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[5\].gen_latches\[2\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[5\]\[2\] net228 dig_ctrl_inst.latch_mem_inst.gclk\[5\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[49\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[49\]\[7\] net189 dig_ctrl_inst.latch_mem_inst.gclk\[49\]
+ sky130_fd_sc_hd__dlxtp_1
X_2500_ VGND VDPWR VDPWR VGND clknet_leaf_5_clk _0097_ net177 net30 sky130_fd_sc_hd__dfrtp_1
X_2431_ VGND VDPWR VDPWR VGND clknet_leaf_13_clk _0039_ net139 dig_ctrl_inst.cpu_inst.data\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_1244_ VGND VDPWR VDPWR VGND _1092_ _1002_ dig_ctrl_inst.spi_addr\[1\] sky130_fd_sc_hd__or2_1
X_2293_ VDPWR VGND VDPWR VGND _0751_ _0920_ _0973_ _0922_ sky130_fd_sc_hd__o21bai_1
X_2362_ VDPWR VGND VDPWR VGND _1039_ dig_ctrl_inst.stb_dd _0999_ _0989_ sky130_fd_sc_hd__a21o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[38\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[38\]\[5\] net204 dig_ctrl_inst.latch_mem_inst.gclk\[38\]
+ sky130_fd_sc_hd__dlxtp_1
X_1313_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[12\] net78 net124
+ net154 sky130_fd_sc_hd__and3_2
XFILLER_0_47_76 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_74_333 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_63_97 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_1175_ VGND VDPWR VDPWR VGND _1020_ _1023_ _1022_ sky130_fd_sc_hd__nand2_1
XANTENNA_23 VGND VDPWR VDPWR VGND _0157_ sky130_fd_sc_hd__diode_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[27\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[27\]\[3\] net217 dig_ctrl_inst.latch_mem_inst.gclk\[27\]
+ sky130_fd_sc_hd__dlxtp_1
XANTENNA_12 VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[56\] sky130_fd_sc_hd__diode_2
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[11\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[11\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[11\] sky130_fd_sc_hd__clkbuf_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[16\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[16\]\[1\] net232 dig_ctrl_inst.latch_mem_inst.gclk\[16\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_65_333 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_25_219 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_17_57 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[9\].gen_latches\[3\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[9\]\[3\] net215 dig_ctrl_inst.latch_mem_inst.gclk\[9\]
+ sky130_fd_sc_hd__dlxtp_1
Xinput10 VGND VDPWR VDPWR VGND net10 ui_in[7] sky130_fd_sc_hd__clkbuf_1
X_1862_ VGND VDPWR VDPWR VGND _0569_ net69 net74 dig_ctrl_inst.latch_mem_inst.RAM\[30\]\[5\]
+ _0159_ dig_ctrl_inst.latch_mem_inst.RAM\[62\]\[5\] sky130_fd_sc_hd__a32o_1
X_1931_ VGND VDPWR VDPWR VGND _0637_ net118 net124 net133 dig_ctrl_inst.latch_mem_inst.RAM\[1\]\[6\]
+ sky130_fd_sc_hd__and4_1
X_1793_ VGND VDPWR VDPWR VGND _0139_ dig_ctrl_inst.latch_mem_inst.RAM\[39\]\[3\] _0499_
+ _0500_ _0501_ _0502_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_3_113 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_58_42 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2414_ VGND VDPWR VDPWR VGND clknet_leaf_13_clk _0022_ net141 dig_ctrl_inst.cpu_inst.ip\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_2345_ VGND VDPWR VDPWR VGND _0095_ net390 _0987_ dig_ctrl_inst.cpu_inst.port_o\[0\]
+ sky130_fd_sc_hd__mux2_1
X_1227_ VDPWR VGND VDPWR VGND _1074_ _1075_ _1067_ _1030_ net293 dig_ctrl_inst.cpu_inst.ip\[0\]
+ sky130_fd_sc_hd__a221oi_4
X_1158_ VDPWR VGND VDPWR VGND _1007_ dig_ctrl_inst.cpu_inst.prev_state\[0\] sky130_fd_sc_hd__inv_2
X_2276_ VGND VDPWR VDPWR VGND _0962_ _0748_ _0956_ _0961_ _0955_ sky130_fd_sc_hd__o211a_1
XFILLER_0_38_333 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_0_127 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_2061_ VGND VDPWR VDPWR VGND net261 _0754_ net257 net288 sky130_fd_sc_hd__or3b_4
X_2130_ VGND VDPWR VDPWR VGND _0258_ _0821_ _0822_ _0257_ sky130_fd_sc_hd__o21ai_1
X_1914_ VGND VDPWR VDPWR VGND _0621_ _0620_ _0603_ _0598_ _0593_ sky130_fd_sc_hd__nor4_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[60\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[60\]\[3\] net223 dig_ctrl_inst.latch_mem_inst.gclk\[60\]
+ sky130_fd_sc_hd__dlxtp_1
X_1845_ VGND VDPWR VDPWR VGND _0553_ net92 net107 net124 dig_ctrl_inst.latch_mem_inst.RAM\[11\]\[4\]
+ sky130_fd_sc_hd__and4_1
X_1776_ VGND VDPWR VDPWR VGND _0120_ dig_ctrl_inst.latch_mem_inst.RAM\[17\]\[3\] _0482_
+ _0483_ _0484_ _0485_ sky130_fd_sc_hd__a2111o_1
X_2328_ VGND VDPWR VDPWR VGND _0080_ dig_ctrl_inst.spi_data_o\[1\] _0180_ dig_ctrl_inst.spi_data_o\[0\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_288 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_2259_ VGND VDPWR VDPWR VGND _0944_ _0946_ _0945_ sky130_fd_sc_hd__nand2_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[25\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[25\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[25\] clknet_leaf_16_clk sky130_fd_sc_hd__dlclkp_1
XFILLER_0_7_260 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1630_ VDPWR VGND VDPWR VGND _0341_ net52 net72 dig_ctrl_inst.latch_mem_inst.RAM\[46\]\[1\]
+ sky130_fd_sc_hd__and3_2
X_1561_ VGND VDPWR VDPWR VGND _0273_ net253 _0274_ sky130_fd_sc_hd__xnor2_1
X_1492_ VGND VDPWR VDPWR VGND _0020_ dig_ctrl_inst.cpu_inst.ip\[1\] _0204_ _0209_
+ sky130_fd_sc_hd__mux2_1
X_2113_ VDPWR VGND VDPWR VGND _0806_ _0755_ _0805_ _0754_ net165 sky130_fd_sc_hd__o2bb2a_1
X_2044_ VGND VDPWR VDPWR VGND _0040_ _0685_ _0741_ net388 sky130_fd_sc_hd__mux2_1
XFILLER_0_44_122 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_188 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_1759_ VDPWR VGND VDPWR VGND _0158_ dig_ctrl_inst.latch_mem_inst.RAM\[9\]\[3\] _1143_
+ _0468_ dig_ctrl_inst.latch_mem_inst.RAM\[61\]\[3\] sky130_fd_sc_hd__a22o_1
X_1828_ VGND VDPWR VDPWR VGND _0536_ net51 net80 net114 dig_ctrl_inst.latch_mem_inst.RAM\[45\]\[4\]
+ sky130_fd_sc_hd__and4_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[53\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[53\]\[2\] net226 dig_ctrl_inst.latch_mem_inst.gclk\[53\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[42\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[42\]\[0\] net243 dig_ctrl_inst.latch_mem_inst.gclk\[42\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_25_57 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[30\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[30\]\[7\] net187 dig_ctrl_inst.latch_mem_inst.gclk\[30\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_41_147 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_1613_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[18\]\[0\] _0121_ _0325_
+ _0151_ dig_ctrl_inst.latch_mem_inst.RAM\[53\]\[0\] _0311_ sky130_fd_sc_hd__a221o_1
X_1544_ VGND VDPWR VDPWR VGND _0254_ _0257_ _0256_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_339 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_26_188 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_1475_ VGND VDPWR VDPWR VGND _0015_ dig_ctrl_inst.cpu_inst.port_o\[4\] _0176_ dig_ctrl_inst.cpu_inst.r0\[4\]
+ sky130_fd_sc_hd__mux2_1
Xfanout219 VGND VDPWR VDPWR VGND net329 net219 sky130_fd_sc_hd__clkbuf_2
Xfanout208 VGND VDPWR VDPWR VGND net209 net208 sky130_fd_sc_hd__clkbuf_2
X_2027_ VDPWR VGND VDPWR VGND _0150_ dig_ctrl_inst.latch_mem_inst.RAM\[21\]\[7\] _0124_
+ _0732_ dig_ctrl_inst.latch_mem_inst.RAM\[52\]\[7\] sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_17_Left_95 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_17_144 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[57\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[57\]\[3\] net220 dig_ctrl_inst.latch_mem_inst.gclk\[57\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_20_309 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
Xdig_ctrl_inst.latch_mem_inst.gen_words\[46\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[46\]\[1\] net234 dig_ctrl_inst.latch_mem_inst.gclk\[46\]
+ sky130_fd_sc_hd__dlxtp_1
X_1191_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.cpu_state\[1\] net248 _1039_
+ _0999_ sky130_fd_sc_hd__nor3_4
X_1260_ VGND VDPWR VDPWR VGND net267 _1108_ dig_ctrl_inst.cpu_inst.r2\[5\] sky130_fd_sc_hd__and2b_1
Xinput8 VGND VDPWR VDPWR VGND net8 ui_in[5] sky130_fd_sc_hd__clkbuf_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[1\].gen_latches\[5\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[1\]\[5\] net202 dig_ctrl_inst.latch_mem_inst.gclk\[1\]
+ sky130_fd_sc_hd__dlxtp_1
X_1527_ VGND VDPWR VDPWR VGND _0240_ _0238_ _0239_ sky130_fd_sc_hd__or2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[23\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[23\]\[6\] net192 dig_ctrl_inst.latch_mem_inst.gclk\[23\]
+ sky130_fd_sc_hd__dlxtp_1
X_1458_ VGND VDPWR VDPWR VGND _0006_ _1096_ _0189_ _0188_ _0184_ sky130_fd_sc_hd__o211a_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[4\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[4\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[4\] clknet_leaf_19_clk sky130_fd_sc_hd__dlclkp_1
X_1389_ VDPWR VGND VDPWR VGND _0150_ net96 net43 sky130_fd_sc_hd__and2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[12\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[12\]\[4\] net214 dig_ctrl_inst.latch_mem_inst.gclk\[12\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[39\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[39\]\[0\] net245 dig_ctrl_inst.latch_mem_inst.gclk\[39\]
+ sky130_fd_sc_hd__dlxtp_1
X_2361_ VGND VDPWR VDPWR VGND _0110_ net353 _0988_ dig_ctrl_inst.cpu_inst.port_o\[7\]
+ sky130_fd_sc_hd__mux2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[5\].gen_latches\[6\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[5\]\[6\] net198 dig_ctrl_inst.latch_mem_inst.gclk\[5\]
+ sky130_fd_sc_hd__dlxtp_1
X_2430_ VGND VDPWR VDPWR VGND clknet_leaf_13_clk _0038_ net139 dig_ctrl_inst.cpu_inst.data\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_2292_ VGND VDPWR VDPWR VGND _0057_ _0972_ _0967_ net359 sky130_fd_sc_hd__mux2_1
X_1243_ VDPWR VGND VDPWR VGND _1091_ _1039_ net162 sky130_fd_sc_hd__and2_1
X_1312_ VDPWR VGND VDPWR VGND _1148_ net125 net79 sky130_fd_sc_hd__and2_1
X_1174_ VGND VDPWR VDPWR VGND net264 _1022_ net265 sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_25_Left_103 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XANTENNA_13 VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[56\] sky130_fd_sc_hd__diode_2
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[50\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[50\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[50\] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_79 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_6_166 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
XANTENNA_24 VGND VDPWR VDPWR VGND _0157_ sky130_fd_sc_hd__diode_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[27\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[27\]\[7\] net189 dig_ctrl_inst.latch_mem_inst.gclk\[27\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_34_Left_112 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_43_Left_121 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[16\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[16\]\[5\] net199 dig_ctrl_inst.latch_mem_inst.gclk\[16\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[32\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[32\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[32\] clknet_leaf_15_clk sky130_fd_sc_hd__dlclkp_1
XPHY_EDGE_ROW_52_Left_130 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_0_309 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_57 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_1930_ VDPWR VGND VDPWR VGND _0636_ net62 net128 dig_ctrl_inst.latch_mem_inst.RAM\[16\]\[6\]
+ sky130_fd_sc_hd__and3_2
X_1792_ VDPWR VGND VDPWR VGND _0501_ net46 net87 dig_ctrl_inst.latch_mem_inst.RAM\[56\]\[3\]
+ sky130_fd_sc_hd__and3_2
Xinput11 VGND VDPWR VDPWR VGND net11 uio_in[0] sky130_fd_sc_hd__clkbuf_1
X_1861_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[11\]\[5\] _1145_ _0568_
+ _0155_ dig_ctrl_inst.latch_mem_inst.RAM\[58\]\[5\] _0567_ sky130_fd_sc_hd__a221o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[9\].gen_latches\[7\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[9\]\[7\] net183 dig_ctrl_inst.latch_mem_inst.gclk\[9\]
+ sky130_fd_sc_hd__dlxtp_1
Xclkbuf_1_0__f_clk VGND VDPWR VDPWR VGND clknet_0_clk clknet_1_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_2344_ VGND VDPWR VDPWR VGND _0802_ _0987_ dig_ctrl_inst.cpu_inst.port_stb_o sky130_fd_sc_hd__nand2_4
X_2413_ VGND VDPWR VDPWR VGND clknet_leaf_9_clk _0021_ net141 dig_ctrl_inst.cpu_inst.ip\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_1226_ VDPWR VGND VDPWR VGND net165 _1039_ net249 _1074_ sky130_fd_sc_hd__a21o_1
X_2275_ VDPWR VGND VDPWR VGND _0956_ _0749_ _0960_ _0961_ sky130_fd_sc_hd__a21oi_1
X_1157_ VDPWR VGND VDPWR VGND _1006_ dig_ctrl_inst.cpu_inst.ip\[5\] sky130_fd_sc_hd__inv_2
XFILLER_0_15_275 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_53_337 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_53_304 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_28_24 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_5_Left_83 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_44_23 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2060_ VGND VDPWR VDPWR VGND net261 net287 _0753_ net257 sky130_fd_sc_hd__nor3b_1
X_1913_ VDPWR VGND VDPWR VGND _0611_ _0619_ _0615_ _0607_ _0620_ sky130_fd_sc_hd__or4_1
X_1844_ VDPWR VGND VDPWR VGND _0552_ net78 net124 dig_ctrl_inst.latch_mem_inst.RAM\[12\]\[4\]
+ sky130_fd_sc_hd__and3_2
X_1775_ VGND VDPWR VDPWR VGND _0484_ net46 net117 net133 dig_ctrl_inst.latch_mem_inst.RAM\[49\]\[3\]
+ sky130_fd_sc_hd__and4_1
X_2327_ VGND VDPWR VDPWR VGND _0079_ dig_ctrl_inst.spi_data_o\[0\] _0180_ net345 sky130_fd_sc_hd__mux2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[60\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[60\]\[7\] net188 dig_ctrl_inst.latch_mem_inst.gclk\[60\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_33_3 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2258_ VGND VDPWR VDPWR VGND _0945_ _0227_ _0921_ sky130_fd_sc_hd__or2_1
X_1209_ VGND VDPWR VDPWR VGND net268 _1057_ dig_ctrl_inst.cpu_inst.r2\[2\] sky130_fd_sc_hd__and2b_1
X_2189_ VGND VDPWR VDPWR VGND _0879_ net162 net165 net166 _1045_ sky130_fd_sc_hd__a31o_1
XFILLER_0_7_294 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_38_131 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_1560_ VGND VDPWR VDPWR VGND _0272_ _0262_ _0273_ _0268_ sky130_fd_sc_hd__o21ai_1
X_2112_ VDPWR VGND VDPWR VGND dig_ctrl_inst.synchronizer_port_i_inst\[0\].out _0802_
+ _0805_ _0804_ dig_ctrl_inst.spi_data_o\[0\] _0803_ sky130_fd_sc_hd__a221o_1
X_1491_ VGND VDPWR VDPWR VGND _0209_ _0208_ _0174_ _0207_ sky130_fd_sc_hd__mux2_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[43\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[43\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[43\] sky130_fd_sc_hd__clkbuf_4
X_2043_ VGND VDPWR VDPWR VGND _0039_ _0622_ _0741_ dig_ctrl_inst.cpu_inst.data\[5\]
+ sky130_fd_sc_hd__mux2_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[9\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[9\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[9\] clknet_leaf_15_clk sky130_fd_sc_hd__dlclkp_1
XFILLER_0_44_134 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_17_337 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_29_197 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1827_ VGND VDPWR VDPWR VGND _0535_ net42 net80 net114 dig_ctrl_inst.latch_mem_inst.RAM\[61\]\[4\]
+ sky130_fd_sc_hd__and4_1
X_1689_ VDPWR VGND VDPWR VGND _0399_ net49 net74 dig_ctrl_inst.latch_mem_inst.RAM\[62\]\[2\]
+ sky130_fd_sc_hd__and3_2
X_1758_ VDPWR VGND VDPWR VGND _0152_ dig_ctrl_inst.latch_mem_inst.RAM\[52\]\[3\] _0150_
+ _0467_ dig_ctrl_inst.latch_mem_inst.RAM\[54\]\[3\] sky130_fd_sc_hd__a22o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[53\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[53\]\[6\] net194 dig_ctrl_inst.latch_mem_inst.gclk\[53\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[42\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[42\]\[4\] net214 dig_ctrl_inst.latch_mem_inst.gclk\[42\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_50_126 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
Xdig_ctrl_inst.latch_mem_inst.gen_words\[31\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[31\]\[2\] net225 dig_ctrl_inst.latch_mem_inst.gclk\[31\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_26_112 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_1474_ VGND VDPWR VDPWR VGND _0014_ dig_ctrl_inst.cpu_inst.port_o\[3\] _0176_ dig_ctrl_inst.cpu_inst.r0\[3\]
+ sky130_fd_sc_hd__mux2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[20\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[20\]\[0\] net245 dig_ctrl_inst.latch_mem_inst.gclk\[20\]
+ sky130_fd_sc_hd__dlxtp_1
X_1612_ VDPWR VGND VDPWR VGND _0308_ _0323_ _0322_ _0306_ _0324_ sky130_fd_sc_hd__or4_1
Xfanout209 VGND VDPWR VDPWR VGND net323 net209 sky130_fd_sc_hd__clkbuf_2
X_1543_ VGND VDPWR VDPWR VGND _0256_ net163 net161 sky130_fd_sc_hd__or2_1
XFILLER_0_5_57 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_9_323 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2026_ VGND VDPWR VDPWR VGND _0126_ dig_ctrl_inst.latch_mem_inst.RAM\[23\]\[7\] _0688_
+ _0689_ _0704_ _0731_ sky130_fd_sc_hd__a2111o_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[37\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[37\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[37\] clknet_leaf_19_clk sky130_fd_sc_hd__dlclkp_1
XFILLER_0_32_137 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[57\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[57\]\[7\] net186 dig_ctrl_inst.latch_mem_inst.gclk\[57\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[2\].gen_latches\[0\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[2\]\[0\] net245 dig_ctrl_inst.latch_mem_inst.gclk\[2\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[46\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[46\]\[5\] net201 dig_ctrl_inst.latch_mem_inst.gclk\[46\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_31_181 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xinput9 VGND VDPWR VDPWR VGND net9 ui_in[6] sky130_fd_sc_hd__clkbuf_1
X_1190_ VDPWR VGND VDPWR VGND _1038_ _1036_ _1025_ _1010_ sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[35\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[35\]\[3\] net216 dig_ctrl_inst.latch_mem_inst.gclk\[35\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[0\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[0\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[0\] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_52_78 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
Xdig_ctrl_inst.latch_mem_inst.gen_words\[24\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[24\]\[1\] net233 dig_ctrl_inst.latch_mem_inst.gclk\[24\]
+ sky130_fd_sc_hd__dlxtp_1
X_1457_ VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_addr\[0\] _0189_ dig_ctrl_inst.spi_addr\[1\]
+ sky130_fd_sc_hd__nand2_1
X_1526_ VGND VDPWR VDPWR VGND _1118_ net159 _0239_ sky130_fd_sc_hd__nor2_1
X_1388_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[51\] net150 _0149_
+ sky130_fd_sc_hd__and2_1
X_2009_ VDPWR VGND VDPWR VGND _0277_ dig_ctrl_inst.latch_mem_inst.RAM\[31\]\[7\] _0132_
+ _0714_ dig_ctrl_inst.latch_mem_inst.RAM\[4\]\[7\] sky130_fd_sc_hd__a22o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[6\].gen_latches\[1\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[6\]\[1\] net232 dig_ctrl_inst.latch_mem_inst.gclk\[6\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[39\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[39\]\[4\] net213 dig_ctrl_inst.latch_mem_inst.gclk\[39\]
+ sky130_fd_sc_hd__dlxtp_1
X_2360_ VGND VDPWR VDPWR VGND _0109_ net383 _0988_ dig_ctrl_inst.cpu_inst.port_o\[6\]
+ sky130_fd_sc_hd__mux2_1
X_1311_ VDPWR VGND VDPWR VGND _1147_ _1047_ net135 net134 _1077_ _1075_ sky130_fd_sc_hd__o2111a_1
X_2291_ VGND VDPWR VDPWR VGND _0903_ _0900_ _0972_ _0751_ sky130_fd_sc_hd__o21ai_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[36\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[36\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[36\] sky130_fd_sc_hd__clkbuf_4
X_1173_ VGND VDPWR VDPWR VGND _1021_ net263 net267 sky130_fd_sc_hd__nor2_4
XFILLER_0_63_44 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_10_Right_10 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1242_ VGND VDPWR VDPWR VGND _1090_ _1089_ _1088_ _1087_ _1086_ net181 sky130_fd_sc_hd__o41a_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[28\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[28\]\[2\] net230 dig_ctrl_inst.latch_mem_inst.gclk\[28\]
+ sky130_fd_sc_hd__dlxtp_1
XANTENNA_25 VGND VDPWR VDPWR VGND _0187_ sky130_fd_sc_hd__diode_2
XANTENNA_14 VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[6\] sky130_fd_sc_hd__diode_2
X_2489_ VGND VDPWR VDPWR VGND clknet_leaf_4_clk _0088_ net177 dig_ctrl_inst.spi_data_i\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[17\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[17\]\[0\] net243 dig_ctrl_inst.latch_mem_inst.gclk\[17\]
+ sky130_fd_sc_hd__dlxtp_1
X_1509_ VGND VDPWR VDPWR VGND _0223_ dig_ctrl_inst.cpu_inst.data\[5\] _0198_ net160
+ sky130_fd_sc_hd__mux2_1
X_1860_ VDPWR VGND VDPWR VGND _0153_ dig_ctrl_inst.latch_mem_inst.RAM\[25\]\[5\] _0128_
+ _0567_ dig_ctrl_inst.latch_mem_inst.RAM\[55\]\[5\] sky130_fd_sc_hd__a22o_1
Xinput12 VGND VDPWR VDPWR VGND net12 uio_in[1] sky130_fd_sc_hd__clkbuf_1
X_1791_ VDPWR VGND VDPWR VGND _0500_ net56 net98 dig_ctrl_inst.latch_mem_inst.RAM\[36\]\[3\]
+ sky130_fd_sc_hd__and3_2
X_2343_ VGND VDPWR VDPWR VGND _0094_ net351 _0986_ dig_ctrl_inst.cpu_inst.port_o\[7\]
+ sky130_fd_sc_hd__mux2_1
X_2274_ VGND VDPWR VDPWR VGND _0960_ _0792_ _0233_ _0172_ _0959_ sky130_fd_sc_hd__a31o_1
X_2412_ VGND VDPWR VDPWR VGND clknet_leaf_9_clk _0020_ net141 dig_ctrl_inst.cpu_inst.ip\[1\]
+ sky130_fd_sc_hd__dfrtp_2
Xclkbuf_leaf_17_clk VGND VDPWR VDPWR VGND clknet_leaf_17_clk clknet_1_0__leaf_clk
+ sky130_fd_sc_hd__clkbuf_8
X_1156_ VDPWR VGND VDPWR VGND _1005_ dig_ctrl_inst.cpu_inst.ip\[4\] sky130_fd_sc_hd__inv_2
X_1225_ VGND VDPWR VDPWR VGND _1073_ _1072_ _1069_ _1070_ _1071_ net181 sky130_fd_sc_hd__o41a_1
XFILLER_0_62_338 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1989_ VDPWR VGND VDPWR VGND _0694_ net51 net93 dig_ctrl_inst.latch_mem_inst.RAM\[38\]\[7\]
+ sky130_fd_sc_hd__and3_2
XFILLER_0_28_69 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_34 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_60_56 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
Xdig_ctrl_inst.latch_mem_inst.gen_words\[61\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[61\]\[2\] net224 dig_ctrl_inst.latch_mem_inst.gclk\[61\]
+ sky130_fd_sc_hd__dlxtp_1
X_1843_ VDPWR VGND VDPWR VGND _0542_ _0550_ _0546_ _0538_ _0551_ sky130_fd_sc_hd__or4_1
X_1912_ VGND VDPWR VDPWR VGND _1143_ dig_ctrl_inst.latch_mem_inst.RAM\[9\]\[5\] _0616_
+ _0617_ _0618_ _0619_ sky130_fd_sc_hd__a2111o_1
Xclkbuf_leaf_6_clk VGND VDPWR VDPWR VGND clknet_leaf_6_clk clknet_1_1__leaf_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_69_43 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
X_1774_ VGND VDPWR VDPWR VGND _0483_ net56 net81 net117 dig_ctrl_inst.latch_mem_inst.RAM\[45\]\[3\]
+ sky130_fd_sc_hd__and4_1
X_2326_ VGND VDPWR VDPWR VGND _0078_ _0182_ dig_ctrl_inst.spi_receiver_inst.spi_cnt\[2\]
+ net174 _0985_ sky130_fd_sc_hd__a31o_1
X_1208_ VDPWR VGND VDPWR VGND _1056_ dig_ctrl_inst.cpu_inst.r3\[2\] net263 net268
+ sky130_fd_sc_hd__and3_2
XPHY_EDGE_ROW_71_Left_149 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[50\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[50\]\[0\] net246 dig_ctrl_inst.latch_mem_inst.gclk\[50\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_26_3 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2257_ VGND VDPWR VDPWR VGND net138 _0944_ _0921_ sky130_fd_sc_hd__nand2_1
X_2188_ VGND VDPWR VDPWR VGND _0878_ net162 net165 net166 _1045_ sky130_fd_sc_hd__and4_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[44\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[44\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[44\] clknet_leaf_19_clk sky130_fd_sc_hd__dlclkp_1
XFILLER_0_53_124 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_53_113 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_39_57 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[29\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[29\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[29\] sky130_fd_sc_hd__clkbuf_4
X_1490_ VDPWR VGND VDPWR VGND dig_ctrl_inst.cpu_inst.ip\[0\] _0208_ dig_ctrl_inst.cpu_inst.ip\[1\]
+ sky130_fd_sc_hd__xor2_1
X_2111_ VGND VDPWR VDPWR VGND _0799_ dig_ctrl_inst.cpu_inst.data\[1\] _0801_ _0804_
+ dig_ctrl_inst.cpu_inst.data\[0\] sky130_fd_sc_hd__and4bb_4
X_2042_ VGND VDPWR VDPWR VGND _0038_ _0565_ _0741_ dig_ctrl_inst.cpu_inst.data\[4\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_88 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_71_66 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_8_Right_8 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1826_ VDPWR VGND VDPWR VGND _0533_ _0529_ _0527_ _0523_ _0534_ sky130_fd_sc_hd__or4_4
XPHY_EDGE_ROW_39_Right_39 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1688_ VGND VDPWR VDPWR VGND _0027_ _0398_ _0276_ net263 sky130_fd_sc_hd__mux2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[54\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[54\]\[1\] net237 dig_ctrl_inst.latch_mem_inst.gclk\[54\]
+ sky130_fd_sc_hd__dlxtp_1
X_1757_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[25\]\[3\] _0128_ _0466_
+ _0151_ dig_ctrl_inst.latch_mem_inst.RAM\[53\]\[3\] _0465_ sky130_fd_sc_hd__a221o_1
X_2309_ VGND VDPWR VDPWR VGND _0069_ _0968_ _0977_ net360 sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_48_Right_48 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_0_91 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_57_Right_57 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_50_116 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_66_Right_66 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1611_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[11\]\[0\] _1145_ _0323_
+ _0117_ dig_ctrl_inst.latch_mem_inst.RAM\[15\]\[0\] _0309_ sky130_fd_sc_hd__a221o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[31\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[31\]\[6\] net191 dig_ctrl_inst.latch_mem_inst.gclk\[31\]
+ sky130_fd_sc_hd__dlxtp_1
X_1473_ VGND VDPWR VDPWR VGND _0013_ dig_ctrl_inst.cpu_inst.port_o\[2\] _0176_ dig_ctrl_inst.cpu_inst.r0\[2\]
+ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_75_Right_75 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1542_ VGND VDPWR VDPWR VGND net163 net161 _0255_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_66 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[20\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[20\]\[4\] net212 dig_ctrl_inst.latch_mem_inst.gclk\[20\]
+ sky130_fd_sc_hd__dlxtp_1
X_2025_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[9\]\[7\] _1143_ _0730_
+ _0135_ dig_ctrl_inst.latch_mem_inst.RAM\[33\]\[7\] _0699_ sky130_fd_sc_hd__a221o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[58\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[58\]\[2\] net229 dig_ctrl_inst.latch_mem_inst.gclk\[58\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_9_313 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1809_ VGND VDPWR VDPWR VGND _1139_ dig_ctrl_inst.latch_mem_inst.RAM\[7\]\[4\] _0514_
+ _0515_ _0516_ _0517_ sky130_fd_sc_hd__a2111o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[47\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[47\]\[0\] net242 dig_ctrl_inst.latch_mem_inst.gclk\[47\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[2\].gen_latches\[4\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[2\]\[4\] net210 dig_ctrl_inst.latch_mem_inst.gclk\[2\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[35\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[35\]\[7\] net184 dig_ctrl_inst.latch_mem_inst.gclk\[35\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_6_305 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[24\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[24\]\[5\] net203 dig_ctrl_inst.latch_mem_inst.gclk\[24\]
+ sky130_fd_sc_hd__dlxtp_1
X_1456_ VDPWR VGND VDPWR VGND _0185_ dig_ctrl_inst.spi_addr\[0\] dig_ctrl_inst.spi_addr\[1\]
+ _0188_ sky130_fd_sc_hd__a21o_1
X_1525_ VDPWR VGND VDPWR VGND _0238_ _1118_ net159 sky130_fd_sc_hd__and2_1
X_1387_ VDPWR VGND VDPWR VGND _0149_ net43 net102 net131 sky130_fd_sc_hd__and3_2
X_2008_ VDPWR VGND VDPWR VGND _0136_ dig_ctrl_inst.latch_mem_inst.RAM\[20\]\[7\] _0123_
+ _0713_ dig_ctrl_inst.latch_mem_inst.RAM\[34\]\[7\] sky130_fd_sc_hd__a22o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[13\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[13\]\[3\] net217 dig_ctrl_inst.latch_mem_inst.gclk\[13\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_9_165 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[6\].gen_latches\[5\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[6\]\[5\] net204 dig_ctrl_inst.latch_mem_inst.gclk\[6\]
+ sky130_fd_sc_hd__dlxtp_1
X_1310_ VGND VDPWR VDPWR VGND _1047_ _1146_ net135 sky130_fd_sc_hd__and2_4
X_2290_ VGND VDPWR VDPWR VGND _0056_ _0971_ _0967_ net375 sky130_fd_sc_hd__mux2_1
X_1241_ VDPWR VGND VDPWR VGND net262 dig_ctrl_inst.cpu_inst.r0\[1\] net266 _1089_
+ sky130_fd_sc_hd__or3_1
X_1172_ VGND VDPWR VDPWR VGND net286 _1019_ _1020_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_15 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_15 VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_data_i\[1\] sky130_fd_sc_hd__diode_2
XANTENNA_26 VGND VDPWR VDPWR VGND _1039_ sky130_fd_sc_hd__diode_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[28\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[28\]\[6\] net194 dig_ctrl_inst.latch_mem_inst.gclk\[28\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_56_3 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_2488_ VGND VDPWR VDPWR VGND clknet_leaf_5_clk _0087_ net177 dig_ctrl_inst.spi_data_i\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_1439_ VDPWR VGND VDPWR VGND _0000_ _0176_ sky130_fd_sc_hd__inv_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[17\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[17\]\[4\] net211 dig_ctrl_inst.latch_mem_inst.gclk\[17\]
+ sky130_fd_sc_hd__dlxtp_1
X_1508_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.ip\[4\] _0220_ _0204_ _0222_
+ _0023_ sky130_fd_sc_hd__a2bb2o_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[49\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[49\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[49\] clknet_leaf_19_clk sky130_fd_sc_hd__dlclkp_1
Xinput13 VGND VDPWR VDPWR VGND net13 uio_in[3] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_141 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1790_ VGND VDPWR VDPWR VGND _0499_ net56 net100 net117 dig_ctrl_inst.latch_mem_inst.RAM\[37\]\[3\]
+ sky130_fd_sc_hd__and4_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[51\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[51\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[51\] clknet_leaf_13_clk sky130_fd_sc_hd__dlclkp_1
X_2411_ VGND VDPWR VDPWR VGND clknet_leaf_13_clk _0019_ net139 dig_ctrl_inst.cpu_inst.ip\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_2342_ VGND VDPWR VDPWR VGND _0093_ net350 _0986_ dig_ctrl_inst.cpu_inst.port_o\[6\]
+ sky130_fd_sc_hd__mux2_1
X_2273_ VDPWR VGND VDPWR VGND dig_ctrl_inst.cpu_inst.data\[7\] _0743_ _0959_ _0825_
+ net138 _0958_ sky130_fd_sc_hd__a221o_1
X_1224_ VDPWR VGND VDPWR VGND net265 net262 dig_ctrl_inst.cpu_inst.r0\[0\] _1072_
+ sky130_fd_sc_hd__or3_1
X_1155_ VDPWR VGND VDPWR VGND _1004_ dig_ctrl_inst.cpu_inst.ip\[3\] sky130_fd_sc_hd__inv_2
X_1988_ VGND VDPWR VDPWR VGND _0693_ net42 net99 net114 dig_ctrl_inst.latch_mem_inst.RAM\[53\]\[7\]
+ sky130_fd_sc_hd__and4_1
Xfanout190 VGND VDPWR VDPWR VGND net328 net190 sky130_fd_sc_hd__clkbuf_2
X_1842_ VGND VDPWR VDPWR VGND _0278_ dig_ctrl_inst.latch_mem_inst.RAM\[5\]\[4\] _0547_
+ _0548_ _0549_ _0550_ sky130_fd_sc_hd__a2111o_1
X_1773_ VGND VDPWR VDPWR VGND _0482_ net66 net91 net104 dig_ctrl_inst.latch_mem_inst.RAM\[27\]\[3\]
+ sky130_fd_sc_hd__and4_1
X_1911_ VGND VDPWR VDPWR VGND _0618_ net52 net80 net115 dig_ctrl_inst.latch_mem_inst.RAM\[45\]\[5\]
+ sky130_fd_sc_hd__and4_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[61\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[61\]\[6\] net191 dig_ctrl_inst.latch_mem_inst.gclk\[61\]
+ sky130_fd_sc_hd__dlxtp_1
X_2325_ VGND VDPWR VDPWR VGND net174 _0985_ dig_ctrl_inst.spi_receiver_inst.stb_o
+ sky130_fd_sc_hd__and2b_1
X_1207_ VDPWR VGND VDPWR VGND _1055_ _1054_ _1025_ _1010_ sky130_fd_sc_hd__and3_2
X_2187_ VDPWR VGND VDPWR VGND _0877_ _0866_ _0876_ sky130_fd_sc_hd__and2_1
X_2256_ VGND VDPWR VDPWR VGND _0943_ _0788_ _0928_ _0932_ _0942_ sky130_fd_sc_hd__o211a_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[50\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[50\]\[4\] net210 dig_ctrl_inst.latch_mem_inst.gclk\[50\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_47_133 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_26_339 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2110_ VGND VDPWR VDPWR VGND _0803_ _0801_ _0800_ dig_ctrl_inst.port_ms_sync_i dig_ctrl_inst.cpu_inst.data\[0\]
+ sky130_fd_sc_hd__and4_1
XFILLER_0_55_57 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
X_2041_ VGND VDPWR VDPWR VGND _0037_ _0505_ _0741_ dig_ctrl_inst.cpu_inst.data\[3\]
+ sky130_fd_sc_hd__mux2_1
X_1825_ VGND VDPWR VDPWR VGND _0128_ dig_ctrl_inst.latch_mem_inst.RAM\[25\]\[4\] _0530_
+ _0531_ _0532_ _0533_ sky130_fd_sc_hd__a2111o_1
X_1756_ VDPWR VGND VDPWR VGND _0465_ net53 net86 dig_ctrl_inst.latch_mem_inst.RAM\[40\]\[3\]
+ sky130_fd_sc_hd__and3_2
X_1687_ VGND VDPWR VDPWR VGND _0397_ _0288_ dig_ctrl_inst.latch_mem_inst.RAM\[0\]\[1\]
+ _0384_ _0398_ sky130_fd_sc_hd__o22a_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[54\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[54\]\[5\] net202 dig_ctrl_inst.latch_mem_inst.gclk\[54\]
+ sky130_fd_sc_hd__dlxtp_1
X_2308_ VGND VDPWR VDPWR VGND _0977_ _0756_ _0175_ net264 net265 sky130_fd_sc_hd__and4_4
X_2239_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.r0\[6\] net41 _0926_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_169 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
Xdig_ctrl_inst.latch_mem_inst.gen_words\[43\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[43\]\[3\] net218 dig_ctrl_inst.latch_mem_inst.gclk\[43\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_23_309 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_8_3 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[32\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[32\]\[1\] net233 dig_ctrl_inst.latch_mem_inst.gclk\[32\]
+ sky130_fd_sc_hd__dlxtp_1
X_1610_ VGND VDPWR VDPWR VGND _0322_ _0310_ _0321_ sky130_fd_sc_hd__or2_1
X_1472_ VGND VDPWR VDPWR VGND _0012_ dig_ctrl_inst.cpu_inst.port_o\[1\] _0176_ dig_ctrl_inst.cpu_inst.r0\[1\]
+ sky130_fd_sc_hd__mux2_1
X_1541_ VGND VDPWR VDPWR VGND net163 _0254_ net161 sky130_fd_sc_hd__nand2_1
X_2024_ VDPWR VGND VDPWR VGND _0722_ _0724_ _0717_ _0729_ sky130_fd_sc_hd__or3_1
X_1808_ VGND VDPWR VDPWR VGND _0516_ net68 _1140_ net108 dig_ctrl_inst.latch_mem_inst.RAM\[27\]\[4\]
+ sky130_fd_sc_hd__and4_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[58\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[58\]\[6\] net198 dig_ctrl_inst.latch_mem_inst.gclk\[58\]
+ sky130_fd_sc_hd__dlxtp_1
X_1739_ VGND VDPWR VDPWR VGND _0435_ _0448_ dig_ctrl_inst.latch_mem_inst.RAM\[0\]\[2\]
+ _0449_ _0434_ _0288_ sky130_fd_sc_hd__o32a_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[47\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[47\]\[4\] net211 dig_ctrl_inst.latch_mem_inst.gclk\[47\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_63_275 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[56\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[56\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[56\] clknet_leaf_0_clk sky130_fd_sc_hd__dlclkp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[36\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[36\]\[2\] net226 dig_ctrl_inst.latch_mem_inst.gclk\[36\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_36_59 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
Xdig_ctrl_inst.latch_mem_inst.gen_words\[25\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[25\]\[0\] net240 dig_ctrl_inst.latch_mem_inst.gclk\[25\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_input_latches\[0\].n_latch VGND VDPWR VDPWR VGND
+ dig_ctrl_inst.latch_mem_inst.wdata\[0\] dig_ctrl_inst.data_out\[0\] clknet_leaf_2_clk
+ sky130_fd_sc_hd__dlxtn_1
XFILLER_0_22_172 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_1524_ VGND VDPWR VDPWR VGND _0230_ _0237_ _0236_ sky130_fd_sc_hd__nand2_1
X_1455_ VDPWR VGND VDPWR VGND _0185_ net382 _0187_ _0005_ sky130_fd_sc_hd__a21oi_1
X_1386_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[50\] net42 net109
+ net148 sky130_fd_sc_hd__and3_2
X_2007_ VDPWR VGND VDPWR VGND _0160_ dig_ctrl_inst.latch_mem_inst.RAM\[57\]\[7\] _0154_
+ _0712_ dig_ctrl_inst.latch_mem_inst.RAM\[63\]\[7\] sky130_fd_sc_hd__a22o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[13\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[13\]\[7\] net183 dig_ctrl_inst.latch_mem_inst.gclk\[13\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[7\].gen_latches\[0\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[7\]\[0\] net247 dig_ctrl_inst.latch_mem_inst.gclk\[7\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_36_253 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[29\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[29\]\[1\] net238 dig_ctrl_inst.latch_mem_inst.gclk\[29\]
+ sky130_fd_sc_hd__dlxtp_1
X_1171_ VGND VDPWR VDPWR VGND net254 net258 _1019_ sky130_fd_sc_hd__or2_4
X_1240_ VGND VDPWR VDPWR VGND net266 _1088_ dig_ctrl_inst.cpu_inst.r2\[1\] sky130_fd_sc_hd__and2b_1
XANTENNA_27 VGND VDPWR VDPWR VGND _1135_ sky130_fd_sc_hd__diode_2
XANTENNA_16 VGND VDPWR VDPWR VGND ui_in[1] sky130_fd_sc_hd__diode_2
XFILLER_0_12_50 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_6_125 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2487_ VGND VDPWR VDPWR VGND clknet_leaf_3_clk net333 net173 dig_ctrl_inst.spi_receiver_inst.spi_sclk_sync
+ sky130_fd_sc_hd__dfrtp_1
X_1507_ VDPWR VGND VDPWR VGND _0222_ _0173_ _0221_ dig_ctrl_inst.cpu_inst.ip\[4\]
+ _0216_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_49_3 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_1369_ VDPWR VGND VDPWR VGND _0141_ net56 net91 net117 sky130_fd_sc_hd__and3_2
X_1438_ VDPWR VGND VDPWR VGND _1020_ _0176_ net266 net264 _0175_ sky130_fd_sc_hd__nand4_4
XFILLER_0_18_275 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_68_175 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xinput14 VGND VDPWR VDPWR VGND net14 uio_in[4] sky130_fd_sc_hd__clkbuf_1
X_2341_ VGND VDPWR VDPWR VGND _0092_ net356 _0986_ dig_ctrl_inst.cpu_inst.port_o\[5\]
+ sky130_fd_sc_hd__mux2_1
X_2410_ VGND VDPWR VDPWR VGND clknet_leaf_6_clk _0018_ net145 dig_ctrl_inst.cpu_inst.port_o\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_1154_ VDPWR VGND VDPWR VGND _1003_ dig_ctrl_inst.spi_addr\[2\] sky130_fd_sc_hd__inv_2
X_2272_ VGND VDPWR VDPWR VGND _0234_ _0785_ _0958_ _0236_ _0957_ _0787_ sky130_fd_sc_hd__o221ai_1
X_1223_ VGND VDPWR VDPWR VGND net262 _1071_ dig_ctrl_inst.cpu_inst.r1\[0\] sky130_fd_sc_hd__and2b_1
XFILLER_0_47_337 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_59_164 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1987_ VGND VDPWR VDPWR VGND _0692_ net51 net102 net131 dig_ctrl_inst.latch_mem_inst.RAM\[35\]\[7\]
+ sky130_fd_sc_hd__and4_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[32\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[32\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[32\] sky130_fd_sc_hd__clkbuf_4
Xfanout180 VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.rst_ni net180 sky130_fd_sc_hd__clkbuf_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[62\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[62\]\[1\] net238 dig_ctrl_inst.latch_mem_inst.gclk\[62\]
+ sky130_fd_sc_hd__dlxtp_1
Xfanout191 VGND VDPWR VDPWR VGND net193 net191 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_60_25 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1910_ VDPWR VGND VDPWR VGND _0617_ net52 net109 dig_ctrl_inst.latch_mem_inst.RAM\[34\]\[5\]
+ sky130_fd_sc_hd__and3_2
XFILLER_0_29_337 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1841_ VDPWR VGND VDPWR VGND _0549_ net97 net123 dig_ctrl_inst.latch_mem_inst.RAM\[4\]\[4\]
+ sky130_fd_sc_hd__and3_2
X_1772_ VGND VDPWR VDPWR VGND _0124_ dig_ctrl_inst.latch_mem_inst.RAM\[21\]\[3\] _0478_
+ _0479_ _0480_ _0481_ sky130_fd_sc_hd__a2111o_1
X_2324_ VGND VDPWR VDPWR VGND _0077_ net355 _0978_ _0984_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_248 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_20_292 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_1206_ VGND VDPWR VDPWR VGND _1054_ _1053_ _1052_ _1051_ _1050_ _1018_ sky130_fd_sc_hd__o41a_4
X_2255_ VDPWR VGND VDPWR VGND _0942_ _0941_ _0936_ _0233_ _0783_ sky130_fd_sc_hd__a211oi_1
X_2186_ VGND VDPWR VDPWR VGND _0876_ _0748_ _0869_ _0875_ _0863_ sky130_fd_sc_hd__o211a_1
XFILLER_0_11_292 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_9_Left_87 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2040_ VGND VDPWR VDPWR VGND _0036_ _0449_ _0741_ dig_ctrl_inst.cpu_inst.data\[2\]
+ sky130_fd_sc_hd__mux2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[55\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[55\]\[0\] net242 dig_ctrl_inst.latch_mem_inst.gclk\[55\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[63\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[63\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[63\] clknet_leaf_18_clk sky130_fd_sc_hd__dlclkp_1
X_1755_ VDPWR VGND VDPWR VGND _0461_ _0463_ _0462_ _0460_ _0464_ sky130_fd_sc_hd__or4_2
X_1686_ VDPWR VGND VDPWR VGND _0386_ _0396_ _0391_ _0287_ _0397_ sky130_fd_sc_hd__or4_1
X_1824_ VGND VDPWR VDPWR VGND _0532_ net54 net100 net117 dig_ctrl_inst.latch_mem_inst.RAM\[37\]\[4\]
+ sky130_fd_sc_hd__and4_1
XFILLER_0_20_61 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2238_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.r0\[5\] _0758_ _0925_ _0050_
+ sky130_fd_sc_hd__o21a_1
X_2307_ VGND VDPWR VDPWR VGND _0068_ _0975_ _0976_ net384 sky130_fd_sc_hd__mux2_1
X_2169_ VGND VDPWR VDPWR VGND _0859_ _0762_ net157 _0761_ sky130_fd_sc_hd__mux2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[43\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[43\]\[7\] net186 dig_ctrl_inst.latch_mem_inst.gclk\[43\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[32\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[32\]\[5\] net201 dig_ctrl_inst.latch_mem_inst.gclk\[32\]
+ sky130_fd_sc_hd__dlxtp_1
X_1540_ VGND VDPWR VDPWR VGND _0248_ _0253_ _0252_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_215 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
Xdig_ctrl_inst.latch_mem_inst.gen_words\[21\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[21\]\[3\] net215 dig_ctrl_inst.latch_mem_inst.gclk\[21\]
+ sky130_fd_sc_hd__dlxtp_1
X_1471_ VGND VDPWR VDPWR VGND _0011_ dig_ctrl_inst.cpu_inst.port_o\[0\] _0176_ dig_ctrl_inst.cpu_inst.r0\[0\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_49 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
X_2023_ VDPWR VGND VDPWR VGND _0711_ _0727_ _0725_ _0710_ _0728_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_59_Left_137 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[59\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[59\]\[1\] net237 dig_ctrl_inst.latch_mem_inst.gclk\[59\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[10\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[10\]\[1\] net235 dig_ctrl_inst.latch_mem_inst.gclk\[10\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[25\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[25\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[25\] sky130_fd_sc_hd__clkbuf_4
X_1807_ VDPWR VGND VDPWR VGND _0515_ net68 net95 dig_ctrl_inst.latch_mem_inst.RAM\[22\]\[4\]
+ sky130_fd_sc_hd__and3_2
XFILLER_0_9_337 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1738_ VDPWR VGND VDPWR VGND _0447_ _0442_ _0439_ _0287_ _0448_ sky130_fd_sc_hd__or4_4
XPHY_EDGE_ROW_68_Left_146 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1669_ VGND VDPWR VDPWR VGND _0151_ dig_ctrl_inst.latch_mem_inst.RAM\[53\]\[1\] _0339_
+ _0340_ _0344_ _0380_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_0_281 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_77_Left_155 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[3\].gen_latches\[3\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[3\]\[3\] net220 dig_ctrl_inst.latch_mem_inst.gclk\[3\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[36\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[36\]\[6\] net195 dig_ctrl_inst.latch_mem_inst.gclk\[36\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_input_latches\[4\].n_latch VDPWR VGND VDPWR VGND
+ dig_ctrl_inst.latch_mem_inst.wdata\[4\] dig_ctrl_inst.data_out\[4\] clknet_leaf_8_clk
+ sky130_fd_sc_hd__dlxtn_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[25\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[25\]\[4\] net208 dig_ctrl_inst.latch_mem_inst.gclk\[25\]
+ sky130_fd_sc_hd__dlxtp_1
X_1454_ VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_addr\[0\] _0186_ _0187_ sky130_fd_sc_hd__nor2_1
X_1523_ VGND VDPWR VDPWR VGND _0236_ _0234_ _0235_ sky130_fd_sc_hd__or2_1
X_1385_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[49\] net156 _0148_
+ sky130_fd_sc_hd__and2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[14\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[14\]\[2\] net228 dig_ctrl_inst.latch_mem_inst.gclk\[14\]
+ sky130_fd_sc_hd__dlxtp_1
X_2006_ VGND VDPWR VDPWR VGND _0709_ _0700_ dig_ctrl_inst.latch_mem_inst.RAM\[10\]\[7\]
+ net123 net294 _0711_ sky130_fd_sc_hd__a311o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[7\].gen_latches\[4\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[7\]\[4\] net212 dig_ctrl_inst.latch_mem_inst.gclk\[7\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_36_287 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_47_15 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_1170_ VGND VDPWR VDPWR VGND _1018_ net254 net258 sky130_fd_sc_hd__nor2_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[29\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[29\]\[5\] net204 dig_ctrl_inst.latch_mem_inst.gclk\[29\]
+ sky130_fd_sc_hd__dlxtp_1
XANTENNA_17 VGND VDPWR VDPWR VGND ui_in[3] sky130_fd_sc_hd__diode_2
XANTENNA_28 VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.port_o\[5\] sky130_fd_sc_hd__diode_2
X_2486_ VGND VDPWR VDPWR VGND clknet_leaf_3_clk net13 net173 dig_ctrl_inst.spi_receiver_inst.synchronizer_spi_sclk.pipe\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[18\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[18\]\[3\] net219 dig_ctrl_inst.latch_mem_inst.gclk\[18\]
+ sky130_fd_sc_hd__dlxtp_1
X_1506_ VGND VDPWR VDPWR VGND _0221_ dig_ctrl_inst.cpu_inst.data\[4\] _0198_ net159
+ sky130_fd_sc_hd__mux2_1
X_1437_ VGND VDPWR VDPWR VGND _0174_ _0175_ dig_ctrl_inst.cpu_inst.skip sky130_fd_sc_hd__nor2_2
X_1299_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[7\] net155 _1139_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_37_70 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1368_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[40\] net53 net86
+ net149 sky130_fd_sc_hd__and3_2
XFILLER_0_18_287 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_17_18 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
Xinput15 VGND VDPWR VDPWR VGND net15 uio_in[5] sky130_fd_sc_hd__buf_1
X_2340_ VGND VDPWR VDPWR VGND _0091_ net348 _0986_ dig_ctrl_inst.cpu_inst.port_o\[4\]
+ sky130_fd_sc_hd__mux2_1
X_2271_ VGND VDPWR VDPWR VGND _0957_ _0791_ _0172_ _0786_ sky130_fd_sc_hd__mux2_1
X_1153_ VDPWR VGND VDPWR VGND _1002_ net251 sky130_fd_sc_hd__inv_2
X_1222_ VGND VDPWR VDPWR VGND net265 _1070_ dig_ctrl_inst.cpu_inst.r2\[0\] sky130_fd_sc_hd__and2b_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[18\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[18\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[18\] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_47_327 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1986_ VDPWR VGND VDPWR VGND _0691_ net48 net78 dig_ctrl_inst.latch_mem_inst.RAM\[60\]\[7\]
+ sky130_fd_sc_hd__and3_2
XFILLER_0_15_246 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_9_clk VGND VDPWR VDPWR VGND clknet_leaf_9_clk clknet_1_1__leaf_clk sky130_fd_sc_hd__clkbuf_8
X_2469_ VGND VDPWR VDPWR VGND clknet_leaf_10_clk _0075_ net142 dig_ctrl_inst.cpu_inst.r3\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_305 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_65_113 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
Xfanout181 VDPWR VGND VDPWR VGND _1021_ net181 sky130_fd_sc_hd__buf_6
Xfanout170 VDPWR VGND VDPWR VGND net170 net171 sky130_fd_sc_hd__buf_2
Xfanout192 VDPWR VGND VDPWR VGND net192 net193 sky130_fd_sc_hd__dlymetal6s2s_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[62\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[62\]\[5\] net205 dig_ctrl_inst.latch_mem_inst.gclk\[62\]
+ sky130_fd_sc_hd__dlxtp_1
X_1840_ VDPWR VGND VDPWR VGND _0548_ net68 net111 dig_ctrl_inst.latch_mem_inst.RAM\[18\]\[4\]
+ sky130_fd_sc_hd__and3_2
XPHY_EDGE_ROW_31_Left_109 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1771_ VGND VDPWR VDPWR VGND _0480_ net62 net80 net103 dig_ctrl_inst.latch_mem_inst.RAM\[31\]\[3\]
+ sky130_fd_sc_hd__and4_1
X_2323_ VGND VDPWR VDPWR VGND _0983_ _0979_ dig_ctrl_inst.spi_receiver_inst.spi_cnt\[2\]
+ _0981_ _0984_ sky130_fd_sc_hd__o22a_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[51\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[51\]\[3\] net222 dig_ctrl_inst.latch_mem_inst.gclk\[51\]
+ sky130_fd_sc_hd__dlxtp_1
X_2254_ VDPWR VGND VDPWR VGND _0938_ _0940_ _0937_ _0941_ sky130_fd_sc_hd__or3_1
X_1205_ VDPWR VGND VDPWR VGND net256 dig_ctrl_inst.cpu_inst.r0\[2\] net260 _1053_
+ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_40_Left_118 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2185_ VDPWR VGND VDPWR VGND _0875_ _0874_ _0871_ _0870_ sky130_fd_sc_hd__and3_2
Xclone18 VGND VDPWR VDPWR VGND net300 _1021_ sky130_fd_sc_hd__clkbuf_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[40\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[40\]\[1\] net234 dig_ctrl_inst.latch_mem_inst.gclk\[40\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_7_287 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1969_ VGND VDPWR VDPWR VGND _0135_ dig_ctrl_inst.latch_mem_inst.RAM\[33\]\[6\] _0632_
+ _0633_ _0639_ _0675_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_11_260 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_135 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
Xdig_ctrl_inst.latch_mem_inst.gen_words\[55\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[55\]\[4\] net208 dig_ctrl_inst.latch_mem_inst.gclk\[55\]
+ sky130_fd_sc_hd__dlxtp_1
X_1823_ VDPWR VGND VDPWR VGND _0531_ net54 net84 dig_ctrl_inst.latch_mem_inst.RAM\[42\]\[4\]
+ sky130_fd_sc_hd__and3_2
Xmax_cap134 VDPWR VGND VDPWR VGND _1094_ net134 sky130_fd_sc_hd__buf_4
X_1754_ VDPWR VGND VDPWR VGND _0129_ dig_ctrl_inst.latch_mem_inst.RAM\[12\]\[3\] _1148_
+ _0463_ dig_ctrl_inst.latch_mem_inst.RAM\[26\]\[3\] sky130_fd_sc_hd__a22o_1
X_1685_ VDPWR VGND VDPWR VGND _0393_ _0395_ _0394_ _0392_ _0396_ sky130_fd_sc_hd__or4_1
X_2237_ VGND VDPWR VDPWR VGND _0920_ _0924_ _0925_ sky130_fd_sc_hd__nand2b_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[44\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[44\]\[2\] net226 dig_ctrl_inst.latch_mem_inst.gclk\[44\]
+ sky130_fd_sc_hd__dlxtp_1
X_2306_ VGND VDPWR VDPWR VGND _0067_ _0974_ _0976_ net363 sky130_fd_sc_hd__mux2_1
X_2168_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.r0\[3\] net41 _0858_ sky130_fd_sc_hd__nor2_1
X_2099_ VGND VDPWR VDPWR VGND _1016_ _0745_ _0792_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_182 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_17_Right_17 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[33\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[33\]\[0\] net240 dig_ctrl_inst.latch_mem_inst.gclk\[33\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_26_Right_26 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_35_Right_35 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1470_ VGND VDPWR VDPWR VGND _0010_ _0196_ dig_ctrl_inst.spi_addr\[5\] _0197_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_1_238 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
Xdig_ctrl_inst.latch_mem_inst.gen_words\[21\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[21\]\[7\] net183 dig_ctrl_inst.latch_mem_inst.gclk\[21\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_44_Right_44 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_5_39 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_53_Right_53 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[59\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[59\]\[5\] net204 dig_ctrl_inst.latch_mem_inst.gclk\[59\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[10\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[10\]\[5\] net204 dig_ctrl_inst.latch_mem_inst.gclk\[10\]
+ sky130_fd_sc_hd__dlxtp_1
X_2022_ VGND VDPWR VDPWR VGND _0727_ _0712_ _0726_ sky130_fd_sc_hd__or2_1
X_1806_ VDPWR VGND VDPWR VGND _0514_ net68 net97 dig_ctrl_inst.latch_mem_inst.RAM\[20\]\[4\]
+ sky130_fd_sc_hd__and3_2
XFILLER_0_25_193 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[48\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[48\]\[3\] net215 dig_ctrl_inst.latch_mem_inst.gclk\[48\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_62_Right_62 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1737_ VDPWR VGND VDPWR VGND _0444_ _0446_ _0445_ _0443_ _0447_ sky130_fd_sc_hd__or4_1
X_1599_ VGND VDPWR VDPWR VGND _0311_ net45 net87 dig_ctrl_inst.latch_mem_inst.RAM\[56\]\[0\]
+ _0146_ dig_ctrl_inst.latch_mem_inst.RAM\[47\]\[0\] sky130_fd_sc_hd__a32o_1
XFILLER_0_0_293 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_1668_ VGND VDPWR VDPWR VGND _0135_ dig_ctrl_inst.latch_mem_inst.RAM\[33\]\[1\] _0352_
+ _0369_ _0372_ _0379_ sky130_fd_sc_hd__a2111o_1
XPHY_EDGE_ROW_71_Right_71 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[3\].gen_latches\[7\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[3\]\[7\] net187 dig_ctrl_inst.latch_mem_inst.gclk\[3\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[37\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[37\]\[1\] net234 dig_ctrl_inst.latch_mem_inst.gclk\[37\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_12_Left_90 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1453_ VDPWR VGND VDPWR VGND _0186_ dig_ctrl_inst.spi_receiver_inst.stb_o dig_ctrl_inst.mode_d
+ net251 sky130_fd_sc_hd__and3_2
XFILLER_0_22_141 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1522_ VDPWR VGND VDPWR VGND _0235_ _0172_ _0233_ sky130_fd_sc_hd__and2_1
X_2005_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[44\]\[7\] _0144_ _0710_
+ _0159_ dig_ctrl_inst.latch_mem_inst.RAM\[62\]\[7\] _0701_ sky130_fd_sc_hd__a221o_1
X_1384_ VDPWR VGND VDPWR VGND _0148_ net50 net118 net132 sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[14\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[14\]\[6\] net192 dig_ctrl_inst.latch_mem_inst.gclk\[14\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_2_29 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_18 VGND VDPWR VDPWR VGND ui_in[7] sky130_fd_sc_hd__diode_2
XANTENNA_29 VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[19\] sky130_fd_sc_hd__diode_2
XFILLER_0_42_247 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1436_ VGND VDPWR VDPWR VGND _0999_ net248 _0174_ dig_ctrl_inst.cpu_inst.cpu_state\[1\]
+ sky130_fd_sc_hd__nand3_2
X_2485_ VGND VDPWR VDPWR VGND clknet_leaf_3_clk net337 net176 dig_ctrl_inst.spi_receiver_inst.spi_cs_sync
+ sky130_fd_sc_hd__dfrtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[18\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[18\]\[7\] net186 dig_ctrl_inst.latch_mem_inst.gclk\[18\]
+ sky130_fd_sc_hd__dlxtp_1
X_1367_ VDPWR VGND VDPWR VGND net86 net53 _0140_ sky130_fd_sc_hd__and2_2
X_1505_ VGND VDPWR VDPWR VGND _0220_ _0204_ _0219_ sky130_fd_sc_hd__or2_1
X_1298_ VDPWR VGND VDPWR VGND _1139_ net101 net106 net126 sky130_fd_sc_hd__and3_2
XFILLER_0_33_236 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_33_225 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[57\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[57\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[57\] sky130_fd_sc_hd__clkbuf_4
X_2270_ VGND VDPWR VDPWR VGND _0933_ _0233_ _0956_ sky130_fd_sc_hd__xnor2_1
X_1221_ VDPWR VGND VDPWR VGND _1069_ dig_ctrl_inst.cpu_inst.r3\[0\] net262 net265
+ sky130_fd_sc_hd__and3_2
X_1152_ VDPWR VGND VDPWR VGND _1001_ dig_ctrl_inst.cpu_inst.ip\[0\] sky130_fd_sc_hd__inv_2
X_1985_ VGND VDPWR VDPWR VGND _0690_ net69 net82 net118 dig_ctrl_inst.latch_mem_inst.RAM\[29\]\[7\]
+ sky130_fd_sc_hd__and4_1
XFILLER_0_23_84 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2399_ VGND VDPWR VDPWR VGND clknet_leaf_3_clk _0008_ net172 dig_ctrl_inst.spi_addr\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_1419_ VDPWR VGND VDPWR VGND _1118_ net249 dig_ctrl_inst.spi_data_o\[4\] dig_ctrl_inst.data_out\[4\]
+ _0162_ sky130_fd_sc_hd__a22o_1
X_2468_ VGND VDPWR VDPWR VGND clknet_leaf_7_clk _0074_ net144 dig_ctrl_inst.cpu_inst.r3\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire40 VGND VDPWR VDPWR VGND net40 _0459_ sky130_fd_sc_hd__clkbuf_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[63\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[63\]\[0\] net242 dig_ctrl_inst.latch_mem_inst.gclk\[63\]
+ sky130_fd_sc_hd__dlxtp_1
Xfanout193 VGND VDPWR VDPWR VGND net194 net193 sky130_fd_sc_hd__clkbuf_2
Xfanout160 VDPWR VGND VDPWR VGND net160 _1110_ sky130_fd_sc_hd__buf_2
Xfanout171 VGND VDPWR VDPWR VGND _1036_ net171 sky130_fd_sc_hd__clkbuf_2
X_1770_ VDPWR VGND VDPWR VGND _0479_ net44 net110 dig_ctrl_inst.latch_mem_inst.RAM\[50\]\[3\]
+ sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[51\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[51\]\[7\] net183 dig_ctrl_inst.latch_mem_inst.gclk\[51\]
+ sky130_fd_sc_hd__dlxtp_1
X_2322_ VGND VDPWR VDPWR VGND _0983_ _0982_ dig_ctrl_inst.spi_receiver_inst.spi_cnt\[1\]
+ dig_ctrl_inst.spi_receiver_inst.spi_cnt\[2\] sky130_fd_sc_hd__a21bo_1
X_1204_ VGND VDPWR VDPWR VGND net256 _1052_ dig_ctrl_inst.cpu_inst.r1\[2\] sky130_fd_sc_hd__and2b_1
X_2253_ VGND VDPWR VDPWR VGND _0787_ _0939_ _0940_ _0230_ sky130_fd_sc_hd__o21ai_1
X_2184_ VDPWR VGND VDPWR VGND _0869_ _0749_ _0873_ _0874_ sky130_fd_sc_hd__a21oi_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[14\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[14\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[14\] clknet_leaf_17_clk sky130_fd_sc_hd__dlclkp_1
X_1899_ VDPWR VGND VDPWR VGND _0606_ net55 net128 dig_ctrl_inst.latch_mem_inst.RAM\[32\]\[5\]
+ sky130_fd_sc_hd__and3_2
X_1968_ VDPWR VGND VDPWR VGND _0664_ _0672_ _0665_ _0673_ _0674_ sky130_fd_sc_hd__or4_4
XFILLER_0_50_71 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
Xdig_ctrl_inst.latch_mem_inst.gen_words\[40\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[40\]\[5\] net202 dig_ctrl_inst.latch_mem_inst.gclk\[40\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_7_266 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_272 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_61_161 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
X_1753_ VDPWR VGND VDPWR VGND _0142_ dig_ctrl_inst.latch_mem_inst.RAM\[15\]\[3\] _0117_
+ _0462_ dig_ctrl_inst.latch_mem_inst.RAM\[42\]\[3\] sky130_fd_sc_hd__a22o_1
X_1822_ VGND VDPWR VDPWR VGND _0530_ net45 net81 net104 dig_ctrl_inst.latch_mem_inst.RAM\[63\]\[4\]
+ sky130_fd_sc_hd__and4_1
X_1684_ VGND VDPWR VDPWR VGND _0141_ dig_ctrl_inst.latch_mem_inst.RAM\[41\]\[1\] _0347_
+ _0351_ _0362_ _0395_ sky130_fd_sc_hd__a2111o_1
X_2167_ VGND VDPWR VDPWR VGND _0047_ _0857_ _0758_ dig_ctrl_inst.cpu_inst.r0\[2\]
+ sky130_fd_sc_hd__mux2_1
X_2236_ VGND VDPWR VDPWR VGND _0923_ _0756_ _0922_ _0754_ _0924_ net41 sky130_fd_sc_hd__o221a_1
X_2305_ VGND VDPWR VDPWR VGND _0066_ _0973_ _0976_ net366 sky130_fd_sc_hd__mux2_1
XFILLER_0_17_3 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[44\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[44\]\[6\] net197 dig_ctrl_inst.latch_mem_inst.gclk\[44\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[0\].gen_latches\[1\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[0\]\[1\] net239 dig_ctrl_inst.latch_mem_inst.gclk\[0\]
+ sky130_fd_sc_hd__dlxtp_1
X_2098_ VGND VDPWR VDPWR VGND _0791_ _1016_ _0744_ sky130_fd_sc_hd__or2_1
XFILLER_0_16_331 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
Xdig_ctrl_inst.latch_mem_inst.gen_words\[33\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[33\]\[4\] net210 dig_ctrl_inst.latch_mem_inst.gclk\[33\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[22\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[22\]\[2\] net226 dig_ctrl_inst.latch_mem_inst.gclk\[22\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[11\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[11\]\[0\] net243 dig_ctrl_inst.latch_mem_inst.gclk\[11\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_66_15 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_2021_ VGND VDPWR VDPWR VGND _0726_ net65 net77 dig_ctrl_inst.latch_mem_inst.RAM\[28\]\[7\]
+ _0127_ dig_ctrl_inst.latch_mem_inst.RAM\[24\]\[7\] sky130_fd_sc_hd__a32o_1
X_1736_ VGND VDPWR VDPWR VGND _0148_ dig_ctrl_inst.latch_mem_inst.RAM\[49\]\[2\] _0400_
+ _0411_ _0413_ _0446_ sky130_fd_sc_hd__a2111o_1
X_1805_ VDPWR VGND VDPWR VGND _0148_ dig_ctrl_inst.latch_mem_inst.RAM\[32\]\[4\] _0134_
+ _0513_ dig_ctrl_inst.latch_mem_inst.RAM\[49\]\[4\] sky130_fd_sc_hd__a22o_1
XFILLER_0_40_153 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1667_ VDPWR VGND VDPWR VGND _1148_ dig_ctrl_inst.latch_mem_inst.RAM\[1\]\[1\] _1130_
+ _0378_ dig_ctrl_inst.latch_mem_inst.RAM\[12\]\[1\] sky130_fd_sc_hd__a22o_1
X_1598_ VDPWR VGND VDPWR VGND _0154_ dig_ctrl_inst.latch_mem_inst.RAM\[22\]\[0\] _0125_
+ _0310_ dig_ctrl_inst.latch_mem_inst.RAM\[57\]\[0\] sky130_fd_sc_hd__a22o_1
XFILLER_0_40_164 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
Xdig_ctrl_inst.latch_mem_inst.gen_words\[48\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[48\]\[7\] net183 dig_ctrl_inst.latch_mem_inst.gclk\[48\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[4\].gen_latches\[2\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[4\]\[2\] net229 dig_ctrl_inst.latch_mem_inst.gclk\[4\]
+ sky130_fd_sc_hd__dlxtp_1
X_2219_ VGND VDPWR VDPWR VGND _0906_ _0244_ _0907_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_48_242 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[37\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[37\]\[5\] net203 dig_ctrl_inst.latch_mem_inst.gclk\[37\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_16_150 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_6_3 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
Xdig_ctrl_inst.latch_mem_inst.gen_words\[26\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[26\]\[3\] net222 dig_ctrl_inst.latch_mem_inst.gclk\[26\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[15\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[15\]\[1\] net235 dig_ctrl_inst.latch_mem_inst.gclk\[15\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_6_309 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1452_ VGND VDPWR VDPWR VGND _1096_ _0185_ _0184_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_337 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1521_ VGND VDPWR VDPWR VGND _0172_ _0233_ _0234_ sky130_fd_sc_hd__nor2_1
X_1383_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[48\] net44 net150
+ net128 sky130_fd_sc_hd__and3_2
X_2004_ VDPWR VGND VDPWR VGND _0138_ dig_ctrl_inst.latch_mem_inst.RAM\[1\]\[7\] _1130_
+ _0709_ dig_ctrl_inst.latch_mem_inst.RAM\[37\]\[7\] sky130_fd_sc_hd__a22o_1
XFILLER_0_9_169 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1719_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[16\]\[2\] _0119_ _0429_
+ _0146_ dig_ctrl_inst.latch_mem_inst.RAM\[47\]\[2\] _0428_ sky130_fd_sc_hd__a221o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[8\].gen_latches\[3\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[8\]\[3\] net217 dig_ctrl_inst.latch_mem_inst.gclk\[8\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[21\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[21\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[21\] sky130_fd_sc_hd__clkbuf_4
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[7\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[7\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[7\] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_337 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[19\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[19\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[19\] clknet_leaf_0_clk sky130_fd_sc_hd__dlclkp_1
XANTENNA_19 VGND VDPWR VDPWR VGND uio_in[0] sky130_fd_sc_hd__diode_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[19\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[19\]\[2\] net229 dig_ctrl_inst.latch_mem_inst.gclk\[19\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_27_201 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_2_312 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_1504_ VDPWR VGND VDPWR VGND _0215_ dig_ctrl_inst.cpu_inst.ip\[4\] _0173_ _0219_
+ sky130_fd_sc_hd__a21oi_1
X_2484_ VGND VDPWR VDPWR VGND clknet_leaf_3_clk net11 net173 dig_ctrl_inst.spi_receiver_inst.synchronizer_spi_cs.pipe\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_1366_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[39\] net156 _0139_
+ sky130_fd_sc_hd__and2_1
X_1435_ VDPWR VGND VDPWR VGND _0173_ _0999_ dig_ctrl_inst.cpu_inst.cpu_state\[1\]
+ net248 sky130_fd_sc_hd__and3_2
X_1297_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[6\] net93 net120
+ net148 sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[21\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[21\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[21\] clknet_leaf_15_clk sky130_fd_sc_hd__dlclkp_1
XFILLER_0_33_19 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1220_ VDPWR VGND VDPWR VGND _1068_ net157 sky130_fd_sc_hd__inv_2
X_1151_ VDPWR VGND VDPWR VGND _1000_ net254 sky130_fd_sc_hd__inv_2
X_1984_ VDPWR VGND VDPWR VGND _0689_ net76 net122 dig_ctrl_inst.latch_mem_inst.RAM\[12\]\[7\]
+ sky130_fd_sc_hd__and3_2
X_2467_ VGND VDPWR VDPWR VGND clknet_leaf_7_clk _0073_ net143 dig_ctrl_inst.cpu_inst.r3\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_2398_ VGND VDPWR VDPWR VGND clknet_leaf_2_clk _0007_ net172 dig_ctrl_inst.spi_addr\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_1418_ VDPWR VGND VDPWR VGND _1036_ net249 dig_ctrl_inst.spi_data_o\[3\] dig_ctrl_inst.data_out\[3\]
+ _0162_ sky130_fd_sc_hd__a22o_1
X_1349_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[30\] net70 net73
+ net153 sky130_fd_sc_hd__and3_2
XFILLER_0_47_3 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
Xfanout172 VGND VDPWR VDPWR VGND net176 net172 sky130_fd_sc_hd__clkbuf_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[63\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[63\]\[4\] net209 dig_ctrl_inst.latch_mem_inst.gclk\[63\]
+ sky130_fd_sc_hd__dlxtp_1
Xfanout183 VGND VDPWR VDPWR VGND net184 net183 sky130_fd_sc_hd__clkbuf_2
Xfanout150 VGND VDPWR VDPWR VGND net151 net150 sky130_fd_sc_hd__clkbuf_2
Xfanout161 VDPWR VGND VDPWR VGND net161 _1090_ sky130_fd_sc_hd__buf_2
Xfanout194 VDPWR VGND VDPWR VGND net194 net322 sky130_fd_sc_hd__buf_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[52\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[52\]\[2\] net225 dig_ctrl_inst.latch_mem_inst.gclk\[52\]
+ sky130_fd_sc_hd__dlxtp_1
X_2321_ VGND VDPWR VDPWR VGND _0982_ dig_ctrl_inst.spi_data_i\[0\] dig_ctrl_inst.spi_receiver_inst.spi_cnt\[0\]
+ dig_ctrl_inst.spi_data_i\[1\] sky130_fd_sc_hd__mux2_1
X_1203_ VDPWR VGND VDPWR VGND _1051_ dig_ctrl_inst.cpu_inst.r3\[2\] net256 net260
+ sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[41\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[41\]\[0\] net240 dig_ctrl_inst.latch_mem_inst.gclk\[41\]
+ sky130_fd_sc_hd__dlxtp_1
X_2252_ VGND VDPWR VDPWR VGND _0939_ _0791_ _0167_ _0786_ sky130_fd_sc_hd__mux2_1
X_2183_ VDPWR VGND VDPWR VGND net159 _0783_ _0873_ _0790_ net170 _0872_ sky130_fd_sc_hd__a221o_1
X_1967_ VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[35\]\[6\] _0137_ _0635_
+ _0642_ _0650_ _0673_ sky130_fd_sc_hd__a2111o_1
X_1898_ VDPWR VGND VDPWR VGND _0605_ net72 net120 dig_ctrl_inst.latch_mem_inst.RAM\[14\]\[5\]
+ sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[14\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[14\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[14\] sky130_fd_sc_hd__clkbuf_4
X_2519_ VDPWR VGND VDPWR VGND uio_oe[0] net269 sky130_fd_sc_hd__buf_2
XFILLER_0_11_251 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[56\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[56\]\[3\] net218 dig_ctrl_inst.latch_mem_inst.gclk\[56\]
+ sky130_fd_sc_hd__dlxtp_1
X_1752_ VGND VDPWR VDPWR VGND _0461_ net69 net79 dig_ctrl_inst.latch_mem_inst.RAM\[28\]\[3\]
+ _0155_ dig_ctrl_inst.latch_mem_inst.RAM\[58\]\[3\] sky130_fd_sc_hd__a32o_1
X_1821_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[40\]\[4\] _0140_ _0529_
+ _0153_ dig_ctrl_inst.latch_mem_inst.RAM\[55\]\[4\] _0528_ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_215 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_10_clk VGND VDPWR VDPWR VGND clknet_leaf_10_clk clknet_1_0__leaf_clk
+ sky130_fd_sc_hd__clkbuf_8
X_1683_ VGND VDPWR VDPWR VGND _1143_ dig_ctrl_inst.latch_mem_inst.RAM\[9\]\[1\] _0349_
+ _0357_ _0361_ _0394_ sky130_fd_sc_hd__a2111o_1
Xmax_cap136 VDPWR VGND VDPWR VGND _1048_ net136 sky130_fd_sc_hd__buf_6
X_2304_ VGND VDPWR VDPWR VGND _0065_ _0972_ _0976_ net378 sky130_fd_sc_hd__mux2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[45\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[45\]\[1\] net234 dig_ctrl_inst.latch_mem_inst.gclk\[45\]
+ sky130_fd_sc_hd__dlxtp_1
X_2235_ VDPWR VGND VDPWR VGND dig_ctrl_inst.spi_data_o\[5\] _0804_ _0923_ dig_ctrl_inst.synchronizer_port_i_inst\[5\].out
+ _0802_ sky130_fd_sc_hd__a22oi_1
X_2166_ VGND VDPWR VDPWR VGND _0756_ _0855_ _0857_ _0754_ _0854_ _0856_ sky130_fd_sc_hd__o221ai_1
X_2097_ VGND VDPWR VDPWR VGND _1016_ _0744_ _0790_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_41 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_3_Right_3 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[0\].gen_latches\[5\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[0\]\[5\] net207 dig_ctrl_inst.latch_mem_inst.gclk\[0\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[0\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[0\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[0\] clknet_leaf_9_clk sky130_fd_sc_hd__dlclkp_1
Xclkbuf_1_1__f_clk VGND VDPWR VDPWR VGND clknet_0_clk clknet_1_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
Xdig_ctrl_inst.latch_mem_inst.gen_words\[22\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[22\]\[6\] net197 dig_ctrl_inst.latch_mem_inst.gclk\[22\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_22_324 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_5_19 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
Xdig_ctrl_inst.latch_mem_inst.gen_words\[11\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[11\]\[4\] net214 dig_ctrl_inst.latch_mem_inst.gclk\[11\]
+ sky130_fd_sc_hd__dlxtp_1
X_2020_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[14\]\[7\] _0116_ _0725_
+ _0140_ dig_ctrl_inst.latch_mem_inst.RAM\[40\]\[7\] _0713_ sky130_fd_sc_hd__a221o_1
XFILLER_0_57_276 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[26\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[26\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[26\] clknet_leaf_0_clk sky130_fd_sc_hd__dlclkp_1
XPHY_EDGE_ROW_28_Left_106 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1735_ VGND VDPWR VDPWR VGND _0114_ dig_ctrl_inst.latch_mem_inst.RAM\[13\]\[2\] _0405_
+ _0414_ _0416_ _0445_ sky130_fd_sc_hd__a2111o_1
X_1804_ VDPWR VGND VDPWR VGND _0149_ dig_ctrl_inst.latch_mem_inst.RAM\[3\]\[4\] _1135_
+ _0512_ dig_ctrl_inst.latch_mem_inst.RAM\[51\]\[4\] sky130_fd_sc_hd__a22o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[49\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[49\]\[2\] net228 dig_ctrl_inst.latch_mem_inst.gclk\[49\]
+ sky130_fd_sc_hd__dlxtp_1
X_1666_ VDPWR VGND VDPWR VGND _0159_ dig_ctrl_inst.latch_mem_inst.RAM\[58\]\[1\] _0155_
+ _0377_ dig_ctrl_inst.latch_mem_inst.RAM\[62\]\[1\] sky130_fd_sc_hd__a22o_1
X_1597_ VGND VDPWR VDPWR VGND _0309_ net57 net95 dig_ctrl_inst.latch_mem_inst.RAM\[38\]\[0\]
+ _0145_ dig_ctrl_inst.latch_mem_inst.RAM\[45\]\[0\] sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_37_Left_115 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[38\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[38\]\[0\] net244 dig_ctrl_inst.latch_mem_inst.gclk\[38\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[4\].gen_latches\[6\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[4\]\[6\] net198 dig_ctrl_inst.latch_mem_inst.gclk\[4\]
+ sky130_fd_sc_hd__dlxtp_1
X_2149_ VGND VDPWR VDPWR VGND _0840_ _0768_ _0780_ sky130_fd_sc_hd__or2_1
X_2218_ VDPWR VGND VDPWR VGND _0240_ _0238_ _0906_ _0884_ sky130_fd_sc_hd__o21bai_1
XPHY_EDGE_ROW_46_Left_124 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_55_Left_133 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[26\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[26\]\[7\] net188 dig_ctrl_inst.latch_mem_inst.gclk\[26\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_64_Left_142 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_73_Left_151 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1520_ VGND VDPWR VDPWR VGND net262 dig_ctrl_inst.cpu_inst.r0\[7\] _0232_ _0233_
+ net265 _0231_ sky130_fd_sc_hd__o32a_4
X_1451_ VGND VDPWR VDPWR VGND _0184_ _1002_ dig_ctrl_inst.mode_d sky130_fd_sc_hd__or2_1
X_1382_ VGND VDPWR VDPWR VGND _1112_ _0147_ _1127_ sky130_fd_sc_hd__and2_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[15\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[15\]\[5\] net199 dig_ctrl_inst.latch_mem_inst.gclk\[15\]
+ sky130_fd_sc_hd__dlxtp_1
X_2003_ VDPWR VGND VDPWR VGND _0708_ net69 net74 dig_ctrl_inst.latch_mem_inst.RAM\[30\]\[7\]
+ sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[60\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[60\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[60\] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_310 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1718_ VDPWR VGND VDPWR VGND _0152_ dig_ctrl_inst.latch_mem_inst.RAM\[2\]\[2\] _1133_
+ _0428_ dig_ctrl_inst.latch_mem_inst.RAM\[54\]\[2\] sky130_fd_sc_hd__a22o_1
XFILLER_0_6_40 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_1649_ VGND VDPWR VDPWR VGND _0360_ net52 net99 net115 dig_ctrl_inst.latch_mem_inst.RAM\[37\]\[1\]
+ sky130_fd_sc_hd__and4_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[8\].gen_latches\[7\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[8\]\[7\] net187 dig_ctrl_inst.latch_mem_inst.gclk\[8\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[19\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[19\]\[6\] net193 dig_ctrl_inst.latch_mem_inst.gclk\[19\]
+ sky130_fd_sc_hd__dlxtp_1
X_2483_ VGND VDPWR VDPWR VGND clknet_leaf_3_clk net336 net173 dig_ctrl_inst.spi_receiver_inst.spi_mosi_sync
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_324 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_1503_ VDPWR VGND VDPWR VGND _0022_ _1004_ _0211_ _0204_ _0218_ sky130_fd_sc_hd__o2bb2a_1
X_1365_ VDPWR VGND VDPWR VGND _0139_ net59 net101 net107 sky130_fd_sc_hd__and3_2
X_1434_ VGND VDPWR VDPWR VGND net27 _1039_ net15 net251 sky130_fd_sc_hd__mux2_1
X_1296_ VDPWR VGND VDPWR VGND _1138_ net136 net135 _1093_ _1077_ _1075_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_68_135 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1150_ VDPWR VGND VDPWR VGND _0999_ dig_ctrl_inst.cpu_inst.cpu_state\[2\] sky130_fd_sc_hd__inv_2
XFILLER_0_23_42 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[5\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[5\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[5\] clknet_leaf_0_clk sky130_fd_sc_hd__dlclkp_1
X_1983_ VDPWR VGND VDPWR VGND _0688_ net47 net110 dig_ctrl_inst.latch_mem_inst.RAM\[50\]\[7\]
+ sky130_fd_sc_hd__and3_2
X_1417_ VDPWR VGND VDPWR VGND _1054_ net250 dig_ctrl_inst.spi_data_o\[2\] dig_ctrl_inst.data_out\[2\]
+ _0162_ sky130_fd_sc_hd__a22o_1
X_2466_ VGND VDPWR VDPWR VGND clknet_leaf_7_clk _0072_ net143 dig_ctrl_inst.cpu_inst.r3\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_2397_ VGND VDPWR VDPWR VGND clknet_leaf_2_clk _0006_ net172 dig_ctrl_inst.spi_addr\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_1279_ VGND VDPWR VDPWR VGND _1120_ _1126_ _1002_ _1127_ _1113_ dig_ctrl_inst.spi_addr\[4\]
+ sky130_fd_sc_hd__o32a_4
X_1348_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[29\] net153 _0131_
+ sky130_fd_sc_hd__and2_1
Xfanout173 VGND VDPWR VDPWR VGND net176 net173 sky130_fd_sc_hd__clkbuf_4
Xfanout162 VGND VDPWR VDPWR VGND net162 _1090_ sky130_fd_sc_hd__buf_1
Xfanout195 VGND VDPWR VDPWR VGND net196 net195 sky130_fd_sc_hd__clkbuf_2
Xfanout151 VGND VDPWR VDPWR VGND net152 net151 sky130_fd_sc_hd__clkbuf_2
Xfanout140 VGND VDPWR VDPWR VGND net147 net140 sky130_fd_sc_hd__clkbuf_4
Xfanout184 VDPWR VGND VDPWR VGND net184 net190 sky130_fd_sc_hd__buf_2
X_2320_ VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_receiver_inst.spi_cnt\[1\] _0981_
+ _0980_ sky130_fd_sc_hd__and2b_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[53\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[53\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[53\] sky130_fd_sc_hd__clkbuf_4
X_2251_ VGND VDPWR VDPWR VGND _0792_ _0228_ _0785_ _0229_ _0938_ sky130_fd_sc_hd__a2bb2o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[52\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[52\]\[6\] net191 dig_ctrl_inst.latch_mem_inst.gclk\[52\]
+ sky130_fd_sc_hd__dlxtp_1
X_1202_ VGND VDPWR VDPWR VGND net256 net260 _1050_ dig_ctrl_inst.cpu_inst.r2\[2\]
+ sky130_fd_sc_hd__and3b_1
X_2182_ VGND VDPWR VDPWR VGND _0825_ net166 _0787_ _0252_ _0872_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_18_97 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1966_ VGND VDPWR VDPWR VGND _1145_ dig_ctrl_inst.latch_mem_inst.RAM\[11\]\[6\] _0637_
+ _0638_ _0649_ _0672_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_34_41 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[41\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[41\]\[4\] net210 dig_ctrl_inst.latch_mem_inst.gclk\[41\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[30\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[30\]\[2\] net230 dig_ctrl_inst.latch_mem_inst.gclk\[30\]
+ sky130_fd_sc_hd__dlxtp_1
X_1897_ VDPWR VGND VDPWR VGND _0604_ net63 net98 dig_ctrl_inst.latch_mem_inst.RAM\[20\]\[5\]
+ sky130_fd_sc_hd__and3_2
X_2449_ VGND VDPWR VDPWR VGND clknet_leaf_6_clk _0057_ net144 dig_ctrl_inst.cpu_inst.r1\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[33\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[33\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[33\] clknet_leaf_12_clk sky130_fd_sc_hd__dlclkp_1
X_2518_ VDPWR VGND VDPWR VGND net16 clknet_leaf_11_clk sky130_fd_sc_hd__buf_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[56\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[56\]\[7\] net188 dig_ctrl_inst.latch_mem_inst.gclk\[56\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_37_160 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1820_ VDPWR VGND VDPWR VGND _0528_ net45 net129 dig_ctrl_inst.latch_mem_inst.RAM\[48\]\[4\]
+ sky130_fd_sc_hd__and3_2
X_1751_ VDPWR VGND VDPWR VGND _0278_ dig_ctrl_inst.latch_mem_inst.RAM\[60\]\[3\] _0157_
+ _0460_ dig_ctrl_inst.latch_mem_inst.RAM\[5\]\[3\] sky130_fd_sc_hd__a22o_1
X_1682_ VGND VDPWR VDPWR VGND _0120_ dig_ctrl_inst.latch_mem_inst.RAM\[17\]\[1\] _0350_
+ _0358_ _0371_ _0393_ sky130_fd_sc_hd__a2111o_1
Xmax_cap137 VGND VDPWR VDPWR VGND _0759_ net137 sky130_fd_sc_hd__clkbuf_2
X_2303_ VGND VDPWR VDPWR VGND _0064_ _0971_ _0976_ net381 sky130_fd_sc_hd__mux2_1
X_2234_ VDPWR VGND VDPWR VGND _1110_ _0922_ _0901_ sky130_fd_sc_hd__xor2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[45\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[45\]\[5\] net199 dig_ctrl_inst.latch_mem_inst.gclk\[45\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[1\].gen_latches\[0\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[1\]\[0\] net240 dig_ctrl_inst.latch_mem_inst.gclk\[1\]
+ sky130_fd_sc_hd__dlxtp_1
X_2165_ VDPWR VGND VDPWR VGND _1060_ _0856_ _0829_ sky130_fd_sc_hd__xor2_1
X_2096_ VGND VDPWR VDPWR VGND _0789_ _0788_ _0787_ _0261_ sky130_fd_sc_hd__a21bo_1
X_1949_ VDPWR VGND VDPWR VGND _0655_ net57 net97 dig_ctrl_inst.latch_mem_inst.RAM\[36\]\[6\]
+ sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[34\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[34\]\[3\] net219 dig_ctrl_inst.latch_mem_inst.gclk\[34\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_0_53 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_0_75 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_43_196 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
X_2522__271 VGND VDPWR VDPWR VGND net271 _2522__271/HI sky130_fd_sc_hd__conb_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[23\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[23\]\[1\] net238 dig_ctrl_inst.latch_mem_inst.gclk\[23\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_13_Right_13 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_22_Right_22 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1803_ VGND VDPWR VDPWR VGND _0511_ _0509_ _0510_ sky130_fd_sc_hd__or2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[5\].gen_latches\[1\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[5\]\[1\] net237 dig_ctrl_inst.latch_mem_inst.gclk\[5\]
+ sky130_fd_sc_hd__dlxtp_1
X_1734_ VDPWR VGND VDPWR VGND _0156_ dig_ctrl_inst.latch_mem_inst.RAM\[26\]\[2\] _0129_
+ _0444_ dig_ctrl_inst.latch_mem_inst.RAM\[59\]\[2\] sky130_fd_sc_hd__a22o_1
X_1596_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[3\]\[0\] _1135_ _0308_
+ _0134_ dig_ctrl_inst.latch_mem_inst.RAM\[32\]\[0\] _0307_ sky130_fd_sc_hd__a221o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[49\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[49\]\[6\] net197 dig_ctrl_inst.latch_mem_inst.gclk\[49\]
+ sky130_fd_sc_hd__dlxtp_1
X_1665_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[54\]\[1\] _0152_ _0376_
+ _0160_ dig_ctrl_inst.latch_mem_inst.RAM\[63\]\[1\] _0375_ sky130_fd_sc_hd__a221o_1
X_2217_ VDPWR VGND VDPWR VGND _0905_ _0900_ _0883_ _0049_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_31_Right_31 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[38\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[38\]\[4\] net213 dig_ctrl_inst.latch_mem_inst.gclk\[38\]
+ sky130_fd_sc_hd__dlxtp_1
X_2148_ VGND VDPWR VDPWR VGND _0777_ _0765_ _0768_ _0763_ _0839_ _0772_ sky130_fd_sc_hd__o221a_1
X_2079_ VGND VDPWR VDPWR VGND net168 _0772_ _0764_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_40_Right_40 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[27\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[27\]\[2\] net227 dig_ctrl_inst.latch_mem_inst.gclk\[27\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[16\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[16\]\[0\] net240 dig_ctrl_inst.latch_mem_inst.gclk\[16\]
+ sky130_fd_sc_hd__dlxtp_1
X_1450_ VDPWR VGND VDPWR VGND net391 _0004_ _0182_ sky130_fd_sc_hd__xor2_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[46\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[46\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[46\] sky130_fd_sc_hd__clkbuf_4
X_1381_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[47\] net152 _0146_
+ sky130_fd_sc_hd__and2_1
X_2002_ VDPWR VGND VDPWR VGND _0707_ net111 net121 dig_ctrl_inst.latch_mem_inst.RAM\[2\]\[7\]
+ sky130_fd_sc_hd__and3_2
XFILLER_0_45_225 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[9\].gen_latches\[2\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[9\]\[2\] net228 dig_ctrl_inst.latch_mem_inst.gclk\[9\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_5_322 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_1717_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[3\]\[2\] _1135_ _0427_
+ _0157_ dig_ctrl_inst.latch_mem_inst.RAM\[60\]\[2\] _0424_ sky130_fd_sc_hd__a221o_1
X_1648_ VDPWR VGND VDPWR VGND _0359_ net52 net86 dig_ctrl_inst.latch_mem_inst.RAM\[40\]\[1\]
+ sky130_fd_sc_hd__and3_2
XFILLER_0_13_155 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1579_ VGND VDPWR VDPWR VGND _0291_ net116 net122 net131 dig_ctrl_inst.latch_mem_inst.RAM\[1\]\[0\]
+ sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_16_Left_94 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_42_228 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2482_ VGND VDPWR VDPWR VGND clknet_leaf_3_clk net12 net173 dig_ctrl_inst.spi_receiver_inst.synchronizer_spi_mosi.pipe\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_1433_ VGND VDPWR VDPWR VGND net26 dig_ctrl_inst.spi_receiver_inst.stb_o net15 dig_ctrl_inst.port_ms_sync_i
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_336 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
X_1502_ VGND VDPWR VDPWR VGND _0174_ _0217_ _0216_ _0218_ sky130_fd_sc_hd__o21a_1
XFILLER_0_10_103 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1295_ VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[5\] _1136_ net118
+ net124 net153 sky130_fd_sc_hd__and4_1
X_1364_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[38\] net51 net93
+ net149 sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[38\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[38\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[38\] clknet_leaf_17_clk sky130_fd_sc_hd__dlclkp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[60\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[60\]\[2\] net224 dig_ctrl_inst.latch_mem_inst.gclk\[60\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_68_125 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_1_Left_79 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[3\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[3\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[3\] sky130_fd_sc_hd__clkbuf_4
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[40\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[40\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[40\] clknet_leaf_17_clk sky130_fd_sc_hd__dlclkp_1
XFILLER_0_59_169 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1982_ VGND VDPWR VDPWR VGND _0687_ net52 net80 net115 dig_ctrl_inst.latch_mem_inst.RAM\[45\]\[7\]
+ sky130_fd_sc_hd__and4_1
X_2465_ VGND VDPWR VDPWR VGND clknet_leaf_8_clk _0071_ net143 dig_ctrl_inst.cpu_inst.r3\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_2396_ VGND VDPWR VDPWR VGND clknet_leaf_3_clk _0005_ net172 dig_ctrl_inst.spi_addr\[0\]
+ sky130_fd_sc_hd__dfrtp_2
X_1416_ VDPWR VGND VDPWR VGND _1084_ net250 dig_ctrl_inst.spi_data_o\[1\] dig_ctrl_inst.data_out\[1\]
+ _0162_ sky130_fd_sc_hd__a22o_1
X_1347_ VDPWR VGND VDPWR VGND _0131_ net70 net82 net118 sky130_fd_sc_hd__and3_2
X_1278_ VDPWR VGND VDPWR VGND _1125_ _1039_ net249 _1126_ sky130_fd_sc_hd__a21o_1
XFILLER_0_64_94 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_42 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_65_106 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_65_139 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_2525__280 VGND VDPWR VDPWR VGND _2525__280/LO net280 sky130_fd_sc_hd__conb_1
Xfanout174 VGND VDPWR VDPWR VGND net176 net174 sky130_fd_sc_hd__clkbuf_4
Xfanout130 VDPWR VGND VDPWR VGND net130 _1095_ sky130_fd_sc_hd__buf_2
Xfanout196 VGND VDPWR VDPWR VGND net196 net198 sky130_fd_sc_hd__buf_1
Xfanout185 VGND VDPWR VDPWR VGND net186 net185 sky130_fd_sc_hd__clkbuf_2
Xfanout163 VGND VDPWR VDPWR VGND _1084_ net163 sky130_fd_sc_hd__buf_8
Xfanout141 VGND VDPWR VDPWR VGND net142 net141 sky130_fd_sc_hd__clkbuf_4
Xfanout152 VGND VDPWR VDPWR VGND _1097_ net152 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_69_Right_69 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[53\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[53\]\[1\] net234 dig_ctrl_inst.latch_mem_inst.gclk\[53\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[39\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[39\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[39\] sky130_fd_sc_hd__clkbuf_4
X_1201_ VGND VDPWR VDPWR VGND _1049_ net182 net297 _1027_ dig_ctrl_inst.cpu_inst.ip\[2\]
+ sky130_fd_sc_hd__o211a_1
X_2250_ VDPWR VGND VDPWR VGND _0825_ dig_ctrl_inst.cpu_inst.data\[6\] _0743_ _0937_
+ net160 sky130_fd_sc_hd__a22o_1
X_2181_ VGND VDPWR VDPWR VGND _0249_ _0786_ net170 _0793_ _0871_ sky130_fd_sc_hd__o22a_1
X_1965_ VDPWR VGND VDPWR VGND _0668_ _0670_ _0669_ _0667_ _0671_ sky130_fd_sc_hd__or4_1
X_2517_ VGND VDPWR VDPWR VGND clknet_leaf_3_clk net251 net173 dig_ctrl_inst.mode_d
+ sky130_fd_sc_hd__dfrtp_1
X_1896_ VDPWR VGND VDPWR VGND _0600_ _0602_ _0601_ _0599_ _0603_ sky130_fd_sc_hd__or4_1
X_2379_ VGND VDPWR VDPWR VGND clknet_leaf_4_clk net339 net174 dig_ctrl_inst.synchronizer_port_i_inst\[7\].out
+ sky130_fd_sc_hd__dfrtp_1
X_2448_ VGND VDPWR VDPWR VGND clknet_leaf_6_clk _0056_ net145 dig_ctrl_inst.cpu_inst.r1\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[30\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[30\]\[6\] net195 dig_ctrl_inst.latch_mem_inst.gclk\[30\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_46_183 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[57\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[57\]\[2\] net224 dig_ctrl_inst.latch_mem_inst.gclk\[57\]
+ sky130_fd_sc_hd__dlxtp_1
X_1750_ VGND VDPWR VDPWR VGND _0459_ _0458_ _0453_ _0451_ _0287_ sky130_fd_sc_hd__nor4_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[46\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[46\]\[0\] net245 dig_ctrl_inst.latch_mem_inst.gclk\[46\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_4_Left_82 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_40_315 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
X_1681_ VGND VDPWR VDPWR VGND _0145_ dig_ctrl_inst.latch_mem_inst.RAM\[45\]\[1\] _0348_
+ _0365_ _0370_ _0392_ sky130_fd_sc_hd__a2111o_1
X_2164_ VDPWR VGND VDPWR VGND dig_ctrl_inst.spi_data_o\[2\] _0804_ _0855_ dig_ctrl_inst.synchronizer_port_i_inst\[2\].out
+ _0802_ sky130_fd_sc_hd__a22oi_1
X_2302_ VGND VDPWR VDPWR VGND _0063_ _0970_ _0976_ net371 sky130_fd_sc_hd__mux2_1
X_2233_ VDPWR VGND VDPWR VGND _0921_ _0878_ _1125_ _1110_ sky130_fd_sc_hd__and3_2
XFILLER_0_29_53 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[1\].gen_latches\[4\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[1\]\[4\] net214 dig_ctrl_inst.latch_mem_inst.gclk\[1\]
+ sky130_fd_sc_hd__dlxtp_1
X_2095_ VGND VDPWR VDPWR VGND _0744_ _1014_ _0788_ sky130_fd_sc_hd__or2_4
X_1948_ VGND VDPWR VDPWR VGND _0654_ net57 _1146_ net107 dig_ctrl_inst.latch_mem_inst.RAM\[47\]\[6\]
+ sky130_fd_sc_hd__and4_1
X_1879_ VGND VDPWR VDPWR VGND _0137_ dig_ctrl_inst.latch_mem_inst.RAM\[35\]\[5\] _0583_
+ _0584_ _0585_ _0586_ sky130_fd_sc_hd__a2111o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[34\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[34\]\[7\] net185 dig_ctrl_inst.latch_mem_inst.gclk\[34\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_31_337 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[10\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[10\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[10\] sky130_fd_sc_hd__clkbuf_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[23\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[23\]\[5\] net201 dig_ctrl_inst.latch_mem_inst.gclk\[23\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[12\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[12\]\[3\] net222 dig_ctrl_inst.latch_mem_inst.gclk\[12\]
+ sky130_fd_sc_hd__dlxtp_1
X_1733_ VDPWR VGND VDPWR VGND _0154_ dig_ctrl_inst.latch_mem_inst.RAM\[25\]\[2\] _0128_
+ _0443_ dig_ctrl_inst.latch_mem_inst.RAM\[57\]\[2\] sky130_fd_sc_hd__a22o_1
X_1802_ VGND VDPWR VDPWR VGND _0510_ net44 net110 dig_ctrl_inst.latch_mem_inst.RAM\[50\]\[4\]
+ _1133_ dig_ctrl_inst.latch_mem_inst.RAM\[2\]\[4\] sky130_fd_sc_hd__a32o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[5\].gen_latches\[5\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[5\]\[5\] net205 dig_ctrl_inst.latch_mem_inst.gclk\[5\]
+ sky130_fd_sc_hd__dlxtp_1
X_1595_ VDPWR VGND VDPWR VGND _0156_ dig_ctrl_inst.latch_mem_inst.RAM\[40\]\[0\] _0140_
+ _0307_ dig_ctrl_inst.latch_mem_inst.RAM\[59\]\[0\] sky130_fd_sc_hd__a22o_1
X_1664_ VGND VDPWR VDPWR VGND _0375_ net50 net88 dig_ctrl_inst.latch_mem_inst.RAM\[56\]\[1\]
+ _0131_ dig_ctrl_inst.latch_mem_inst.RAM\[29\]\[1\] sky130_fd_sc_hd__a32o_1
XFILLER_0_13_337 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_0_253 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_2216_ VGND VDPWR VDPWR VGND _0904_ _0756_ _0903_ _0754_ _0905_ net41 sky130_fd_sc_hd__o221a_1
X_2147_ VDPWR VGND VDPWR VGND _0838_ _0264_ _0760_ _0836_ _0770_ _0837_ sky130_fd_sc_hd__o32a_1
X_2078_ VDPWR VGND VDPWR VGND _0760_ _0770_ _0264_ _0771_ sky130_fd_sc_hd__or3_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[45\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[45\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[45\] clknet_leaf_16_clk sky130_fd_sc_hd__dlclkp_1
XFILLER_0_31_134 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
Xdig_ctrl_inst.latch_mem_inst.gen_words\[27\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[27\]\[6\] net198 dig_ctrl_inst.latch_mem_inst.gclk\[27\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[16\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[16\]\[4\] net208 dig_ctrl_inst.latch_mem_inst.gclk\[16\]
+ sky130_fd_sc_hd__dlxtp_1
X_1380_ VGND VDPWR VDPWR VGND _0146_ net104 net81 net54 sky130_fd_sc_hd__and3_4
X_2001_ VGND VDPWR VDPWR VGND _0706_ net42 net80 net115 dig_ctrl_inst.latch_mem_inst.RAM\[61\]\[7\]
+ sky130_fd_sc_hd__and4_1
XFILLER_0_42_75 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
Xdig_ctrl_inst.latch_mem_inst.gen_words\[9\].gen_latches\[6\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[9\]\[6\] net197 dig_ctrl_inst.latch_mem_inst.gclk\[9\]
+ sky130_fd_sc_hd__dlxtp_1
X_1716_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[35\]\[2\] _0137_ _0426_
+ _0145_ dig_ctrl_inst.latch_mem_inst.RAM\[45\]\[2\] _0425_ sky130_fd_sc_hd__a221o_1
X_1578_ VGND VDPWR VDPWR VGND _0290_ net71 net101 net108 dig_ctrl_inst.latch_mem_inst.RAM\[23\]\[0\]
+ sky130_fd_sc_hd__and4_1
X_1647_ VGND VDPWR VDPWR VGND _0358_ net66 net105 net133 dig_ctrl_inst.latch_mem_inst.RAM\[19\]\[1\]
+ sky130_fd_sc_hd__and4_1
Xrebuffer20 VDPWR VGND VDPWR VGND net302 net303 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_4_3 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_2481_ VDPWR VGND VDPWR VGND clknet_leaf_3_clk net344 dig_ctrl_inst.spi_receiver_inst.spi_sclk_delayed
+ sky130_fd_sc_hd__dfxtp_1
X_1432_ VDPWR VGND VDPWR VGND _0162_ net250 dig_ctrl_inst.spi_data_o\[7\] dig_ctrl_inst.data_out\[7\]
+ _0172_ sky130_fd_sc_hd__a22o_1
X_1363_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[37\] net156 _0138_
+ sky130_fd_sc_hd__and2_1
X_1501_ VGND VDPWR VDPWR VGND _0217_ dig_ctrl_inst.cpu_inst.data\[3\] _0198_ net169
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_148 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1294_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[4\] net97 net125
+ net154 sky130_fd_sc_hd__and3_2
XFILLER_0_53_41 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[60\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[60\]\[6\] net322 dig_ctrl_inst.latch_mem_inst.gclk\[60\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_17_281 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_1981_ VGND VDPWR VDPWR VGND _0686_ dig_ctrl_inst.latch_mem_inst.RAM\[0\]\[7\] _0288_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_15_229 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
X_2395_ VGND VDPWR VDPWR VGND clknet_leaf_6_clk net340 net180 dig_ctrl_inst.port_ms_sync_i
+ sky130_fd_sc_hd__dfrtp_1
X_1415_ VDPWR VGND VDPWR VGND _1067_ net250 dig_ctrl_inst.spi_data_o\[0\] dig_ctrl_inst.data_out\[0\]
+ _0162_ sky130_fd_sc_hd__a22o_1
X_1346_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[28\] net70 net78
+ net153 sky130_fd_sc_hd__and3_2
X_2464_ VGND VDPWR VDPWR VGND clknet_leaf_10_clk _0070_ net139 dig_ctrl_inst.cpu_inst.r3\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_1277_ VGND VDPWR VDPWR VGND _1021_ _1121_ _1122_ _1123_ _1124_ _1125_ sky130_fd_sc_hd__o41a_2
XFILLER_0_14_273 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
Xfanout120 VDPWR VGND VDPWR VGND net120 net122 sky130_fd_sc_hd__buf_2
Xfanout131 VDPWR VGND VDPWR VGND net131 net133 sky130_fd_sc_hd__buf_2
Xfanout142 VDPWR VGND VDPWR VGND net142 net147 sky130_fd_sc_hd__buf_2
Xfanout175 VGND VDPWR VDPWR VGND net176 net175 sky130_fd_sc_hd__clkbuf_2
Xfanout153 VGND VDPWR VDPWR VGND net154 net153 sky130_fd_sc_hd__clkbuf_2
Xfanout186 VGND VDPWR VDPWR VGND net190 net186 sky130_fd_sc_hd__clkbuf_2
Xfanout197 VGND VDPWR VDPWR VGND net198 net197 sky130_fd_sc_hd__clkbuf_2
Xfanout164 VDPWR VGND VDPWR VGND net164 net295 sky130_fd_sc_hd__buf_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[53\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[53\]\[5\] net199 dig_ctrl_inst.latch_mem_inst.gclk\[53\]
+ sky130_fd_sc_hd__dlxtp_1
X_1200_ VGND VDPWR VDPWR VGND _1008_ _1048_ _1038_ net249 _1029_ _1046_ sky130_fd_sc_hd__o41ai_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[42\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[42\]\[3\] net222 dig_ctrl_inst.latch_mem_inst.gclk\[42\]
+ sky130_fd_sc_hd__dlxtp_1
X_2180_ VDPWR VGND VDPWR VGND _0870_ dig_ctrl_inst.cpu_inst.data\[3\] _0743_ _0250_
+ _0785_ sky130_fd_sc_hd__o2bb2a_1
X_1964_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[29\]\[6\] _0131_ _0670_
+ _0144_ dig_ctrl_inst.latch_mem_inst.RAM\[44\]\[6\] _0662_ sky130_fd_sc_hd__a221o_1
X_1895_ VDPWR VGND VDPWR VGND _0160_ dig_ctrl_inst.latch_mem_inst.RAM\[47\]\[5\] _0146_
+ _0602_ dig_ctrl_inst.latch_mem_inst.RAM\[63\]\[5\] sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_13_clk VGND VDPWR VDPWR VGND clknet_leaf_13_clk clknet_1_0__leaf_clk
+ sky130_fd_sc_hd__clkbuf_8
Xdig_ctrl_inst.latch_mem_inst.gen_words\[31\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[31\]\[1\] net233 dig_ctrl_inst.latch_mem_inst.gclk\[31\]
+ sky130_fd_sc_hd__dlxtp_1
X_2447_ VGND VDPWR VDPWR VGND clknet_leaf_8_clk _0055_ net146 dig_ctrl_inst.cpu_inst.r1\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_2516_ VGND VDPWR VDPWR VGND clknet_leaf_8_clk _0113_ net143 dig_ctrl_inst.cpu_inst.cpu_state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_2378_ VGND VDPWR VDPWR VGND clknet_leaf_3_clk net10 net173 dig_ctrl_inst.synchronizer_port_i_inst\[7\].pipe\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_1329_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[19\] net154 _0122_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_45_3 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[57\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[57\]\[6\] net194 dig_ctrl_inst.latch_mem_inst.gclk\[57\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[52\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[52\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[52\] clknet_leaf_12_clk sky130_fd_sc_hd__dlclkp_1
X_1680_ VDPWR VGND VDPWR VGND _0388_ _0390_ _0389_ _0387_ _0391_ sky130_fd_sc_hd__or4_1
X_2301_ VGND VDPWR VDPWR VGND _0062_ _0969_ _0976_ net362 sky130_fd_sc_hd__mux2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[46\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[46\]\[4\] net210 dig_ctrl_inst.latch_mem_inst.gclk\[46\]
+ sky130_fd_sc_hd__dlxtp_1
Xclkbuf_leaf_2_clk VGND VDPWR VDPWR VGND clknet_leaf_2_clk clknet_1_1__leaf_clk sky130_fd_sc_hd__clkbuf_8
X_2232_ VGND VDPWR VDPWR VGND _0920_ _0910_ _0907_ _0788_ _0919_ sky130_fd_sc_hd__o211ai_2
X_2163_ VGND VDPWR VDPWR VGND _0854_ _0788_ _0853_ _0851_ _0841_ sky130_fd_sc_hd__o211a_1
X_2094_ VDPWR VGND VDPWR VGND _0787_ _0742_ _0745_ sky130_fd_sc_hd__or2_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[35\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[35\]\[2\] net224 dig_ctrl_inst.latch_mem_inst.gclk\[35\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_9_53 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_16_302 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1947_ VDPWR VGND VDPWR VGND _0653_ net75 net120 dig_ctrl_inst.latch_mem_inst.RAM\[14\]\[6\]
+ sky130_fd_sc_hd__and3_2
X_1878_ VGND VDPWR VDPWR VGND _0585_ net62 net81 net102 dig_ctrl_inst.latch_mem_inst.RAM\[31\]\[5\]
+ sky130_fd_sc_hd__and4_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[24\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[24\]\[0\] net240 dig_ctrl_inst.latch_mem_inst.gclk\[24\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_19_140 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[12\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[12\]\[7\] net183 dig_ctrl_inst.latch_mem_inst.gclk\[12\]
+ sky130_fd_sc_hd__dlxtp_1
X_1732_ VGND VDPWR VDPWR VGND _0442_ _0440_ _0441_ sky130_fd_sc_hd__or2_1
X_1663_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[4\]\[1\] _0277_ _0374_
+ _0278_ dig_ctrl_inst.latch_mem_inst.RAM\[5\]\[1\] _0373_ sky130_fd_sc_hd__a221o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[6\].gen_latches\[0\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[6\]\[0\] net241 dig_ctrl_inst.latch_mem_inst.gclk\[6\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_13_316 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_1801_ VGND VDPWR VDPWR VGND _0509_ net55 net75 dig_ctrl_inst.latch_mem_inst.RAM\[46\]\[4\]
+ _0137_ dig_ctrl_inst.latch_mem_inst.RAM\[35\]\[4\] sky130_fd_sc_hd__a32o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[39\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[39\]\[3\] net218 dig_ctrl_inst.latch_mem_inst.gclk\[39\]
+ sky130_fd_sc_hd__dlxtp_1
X_1594_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[2\]\[0\] _1133_ _0306_
+ _0139_ dig_ctrl_inst.latch_mem_inst.RAM\[39\]\[0\] _0305_ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_265 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Right_7 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2215_ VDPWR VGND VDPWR VGND dig_ctrl_inst.spi_data_o\[4\] _0804_ _0904_ dig_ctrl_inst.synchronizer_port_i_inst\[4\].out
+ _0802_ sky130_fd_sc_hd__a22oi_1
X_2077_ VGND VDPWR VDPWR VGND net163 _0770_ _0769_ sky130_fd_sc_hd__nand2b_2
X_2146_ VGND VDPWR VDPWR VGND _0837_ _0766_ net157 _0762_ sky130_fd_sc_hd__mux2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[28\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[28\]\[1\] net236 dig_ctrl_inst.latch_mem_inst.gclk\[28\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_31_113 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_24_Left_102 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_33_Left_111 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_42_Left_120 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2000_ VGND VDPWR VDPWR VGND _0705_ net51 net90 net114 dig_ctrl_inst.latch_mem_inst.RAM\[41\]\[7\]
+ sky130_fd_sc_hd__and4_1
X_1646_ VGND VDPWR VDPWR VGND _0357_ net61 net90 net115 dig_ctrl_inst.latch_mem_inst.RAM\[25\]\[1\]
+ sky130_fd_sc_hd__and4_1
X_1715_ VDPWR VGND VDPWR VGND _0158_ dig_ctrl_inst.latch_mem_inst.RAM\[32\]\[2\] _0134_
+ _0425_ dig_ctrl_inst.latch_mem_inst.RAM\[61\]\[2\] sky130_fd_sc_hd__a22o_1
X_1577_ VDPWR VGND VDPWR VGND _0289_ net58 net111 dig_ctrl_inst.latch_mem_inst.RAM\[34\]\[0\]
+ sky130_fd_sc_hd__and3_2
XFILLER_0_6_98 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xrebuffer21 VGND VDPWR VDPWR VGND net303 _1076_ sky130_fd_sc_hd__clkbuf_1
Xrebuffer10 VDPWR VGND VDPWR VGND net292 _1026_ sky130_fd_sc_hd__dlygate4sd1_1
X_2129_ VDPWR VGND VDPWR VGND _0258_ _0257_ _0788_ _0821_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_36_249 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2480_ VGND VDPWR VDPWR VGND clknet_leaf_2_clk _0086_ net180 dig_ctrl_inst.spi_data_o\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_230 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1500_ VGND VDPWR VDPWR VGND _0174_ _0216_ _0215_ sky130_fd_sc_hd__nand2_1
X_1293_ VDPWR VGND VDPWR VGND _1137_ net136 net135 net134 _1077_ _1075_ sky130_fd_sc_hd__o2111a_1
X_1362_ VDPWR VGND VDPWR VGND _0138_ net57 net101 net118 sky130_fd_sc_hd__and3_2
X_1431_ VGND VDPWR VDPWR VGND _0172_ _0171_ _0170_ _0169_ _0168_ _1018_ sky130_fd_sc_hd__o41a_4
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[42\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[42\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[42\] sky130_fd_sc_hd__clkbuf_4
X_1629_ VDPWR VGND VDPWR VGND _0340_ net47 net76 dig_ctrl_inst.latch_mem_inst.RAM\[60\]\[1\]
+ sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[61\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[61\]\[1\] net232 dig_ctrl_inst.latch_mem_inst.gclk\[61\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[57\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[57\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[57\] clknet_leaf_16_clk sky130_fd_sc_hd__dlclkp_1
XFILLER_0_17_293 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_17_271 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_59_105 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1980_ VGND VDPWR VDPWR VGND _0032_ _0685_ _0276_ dig_ctrl_inst.cpu_inst.instr\[6\]
+ sky130_fd_sc_hd__mux2_1
X_2532_ VDPWR VGND VDPWR VGND uio_out[5] net278 sky130_fd_sc_hd__buf_2
Xrebuffer1 VDPWR VGND VDPWR VGND _1017_ net283 sky130_fd_sc_hd__buf_6
X_2463_ VGND VDPWR VDPWR VGND clknet_leaf_11_clk _0069_ net140 dig_ctrl_inst.cpu_inst.r3\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_1414_ VGND VDPWR VDPWR VGND _1040_ _0162_ net250 sky130_fd_sc_hd__nor2_2
X_2394_ VGND VDPWR VDPWR VGND clknet_leaf_6_clk net1 net180 dig_ctrl_inst.synchronizer_port_ms_i_inst.pipe\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_1276_ VDPWR VGND VDPWR VGND net263 dig_ctrl_inst.cpu_inst.r0\[4\] net268 _1124_
+ sky130_fd_sc_hd__or3_1
X_1345_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[27\] net155 _0130_
+ sky130_fd_sc_hd__and2_1
Xfanout132 VGND VDPWR VDPWR VGND net133 net132 sky130_fd_sc_hd__clkbuf_4
Xfanout143 VGND VDPWR VDPWR VGND net147 net143 sky130_fd_sc_hd__clkbuf_4
Xfanout154 VGND VDPWR VDPWR VGND net155 net154 sky130_fd_sc_hd__clkbuf_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[54\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[54\]\[0\] net240 dig_ctrl_inst.latch_mem_inst.gclk\[54\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_14_285 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
Xfanout110 VDPWR VGND VDPWR VGND net110 net112 sky130_fd_sc_hd__buf_2
Xfanout121 VGND VDPWR VDPWR VGND net122 net121 sky130_fd_sc_hd__clkbuf_2
Xfanout165 VDPWR VGND VDPWR VGND _1073_ net165 sky130_fd_sc_hd__buf_6
Xfanout176 VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.rst_ni net176 sky130_fd_sc_hd__clkbuf_2
Xfanout187 VDPWR VGND VDPWR VGND net187 net188 sky130_fd_sc_hd__buf_2
Xfanout198 VDPWR VGND VDPWR VGND net198 net322 sky130_fd_sc_hd__buf_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[42\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[42\]\[7\] net188 dig_ctrl_inst.latch_mem_inst.gclk\[42\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_18_23 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1894_ VGND VDPWR VDPWR VGND _0601_ net45 net111 dig_ctrl_inst.latch_mem_inst.RAM\[50\]\[5\]
+ _0138_ dig_ctrl_inst.latch_mem_inst.RAM\[37\]\[5\] sky130_fd_sc_hd__a32o_1
X_1963_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[20\]\[6\] _0123_ _0669_
+ _0278_ dig_ctrl_inst.latch_mem_inst.RAM\[5\]\[6\] _0661_ sky130_fd_sc_hd__a221o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[31\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[31\]\[5\] net199 dig_ctrl_inst.latch_mem_inst.gclk\[31\]
+ sky130_fd_sc_hd__dlxtp_1
X_2515_ VGND VDPWR VDPWR VGND clknet_leaf_9_clk _0112_ net142 dig_ctrl_inst.cpu_inst.cpu_state\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_2446_ VGND VDPWR VDPWR VGND clknet_leaf_9_clk _0054_ net141 dig_ctrl_inst.cpu_inst.r1\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_3 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1259_ VDPWR VGND VDPWR VGND _1107_ dig_ctrl_inst.cpu_inst.r3\[5\] net263 net267
+ sky130_fd_sc_hd__and3_2
X_2377_ VGND VDPWR VDPWR VGND clknet_leaf_4_clk _0004_ net177 dig_ctrl_inst.spi_receiver_inst.spi_cnt\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_1328_ VDPWR VGND VDPWR VGND _0122_ net70 net107 net132 sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[20\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[20\]\[3\] net220 dig_ctrl_inst.latch_mem_inst.gclk\[20\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_19_333 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[58\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[58\]\[1\] net238 dig_ctrl_inst.latch_mem_inst.gclk\[58\]
+ sky130_fd_sc_hd__dlxtp_1
X_2231_ VGND VDPWR VDPWR VGND _0919_ _0750_ _0912_ _0917_ _0918_ sky130_fd_sc_hd__o211a_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[2\].gen_latches\[3\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[2\]\[3\] net215 dig_ctrl_inst.latch_mem_inst.gclk\[2\]
+ sky130_fd_sc_hd__dlxtp_1
X_2300_ VGND VDPWR VDPWR VGND _0061_ _0968_ _0976_ net379 sky130_fd_sc_hd__mux2_1
X_2162_ VGND VDPWR VDPWR VGND _0852_ _0248_ _0853_ sky130_fd_sc_hd__xnor2_1
X_2093_ VGND VDPWR VDPWR VGND net252 _0786_ net253 _0745_ sky130_fd_sc_hd__or3b_4
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[35\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[35\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[35\] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_28_163 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[35\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[35\]\[6\] net194 dig_ctrl_inst.latch_mem_inst.gclk\[35\]
+ sky130_fd_sc_hd__dlxtp_1
X_1946_ VDPWR VGND VDPWR VGND _0652_ net57 net95 dig_ctrl_inst.latch_mem_inst.RAM\[38\]\[6\]
+ sky130_fd_sc_hd__and3_2
XFILLER_0_43_122 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1877_ VGND VDPWR VDPWR VGND _0584_ net44 net99 net114 dig_ctrl_inst.latch_mem_inst.RAM\[53\]\[5\]
+ sky130_fd_sc_hd__and4_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[24\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[24\]\[4\] net211 dig_ctrl_inst.latch_mem_inst.gclk\[24\]
+ sky130_fd_sc_hd__dlxtp_1
X_2429_ VGND VDPWR VDPWR VGND clknet_leaf_9_clk _0037_ net141 dig_ctrl_inst.cpu_inst.data\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[13\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[13\]\[2\] net229 dig_ctrl_inst.latch_mem_inst.gclk\[13\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_34_166 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1800_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[23\]\[4\] _0126_ _0508_
+ _0279_ dig_ctrl_inst.latch_mem_inst.RAM\[6\]\[4\] _0507_ sky130_fd_sc_hd__a221o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[6\].gen_latches\[4\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[6\]\[4\] net211 dig_ctrl_inst.latch_mem_inst.gclk\[6\]
+ sky130_fd_sc_hd__dlxtp_1
Xwire182 VGND VDPWR VDPWR VGND _1009_ net182 sky130_fd_sc_hd__clkbuf_2
X_1662_ VDPWR VGND VDPWR VGND _0148_ dig_ctrl_inst.latch_mem_inst.RAM\[42\]\[1\] _0142_
+ _0373_ dig_ctrl_inst.latch_mem_inst.RAM\[49\]\[1\] sky130_fd_sc_hd__a22o_1
X_1731_ VGND VDPWR VDPWR VGND _0441_ net57 net73 dig_ctrl_inst.latch_mem_inst.RAM\[46\]\[2\]
+ _0138_ dig_ctrl_inst.latch_mem_inst.RAM\[37\]\[2\] sky130_fd_sc_hd__a32o_1
XFILLER_0_13_328 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_2214_ VGND VDPWR VDPWR VGND _0901_ _0903_ _0902_ sky130_fd_sc_hd__nand2_1
X_1593_ VDPWR VGND VDPWR VGND _0143_ dig_ctrl_inst.latch_mem_inst.RAM\[20\]\[0\] _0123_
+ _0305_ dig_ctrl_inst.latch_mem_inst.RAM\[43\]\[0\] sky130_fd_sc_hd__a22o_1
XFILLER_0_0_277 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[39\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[39\]\[7\] net189 dig_ctrl_inst.latch_mem_inst.gclk\[39\]
+ sky130_fd_sc_hd__dlxtp_1
X_2076_ VGND VDPWR VDPWR VGND net253 dig_ctrl_inst.cpu_inst.instr\[6\] dig_ctrl_inst.cpu_inst.instr\[7\]
+ net252 _0769_ sky130_fd_sc_hd__and4bb_1
X_2145_ VGND VDPWR VDPWR VGND _0836_ net163 _0769_ sky130_fd_sc_hd__nand2_2
X_1929_ VDPWR VGND VDPWR VGND _0635_ net64 net86 dig_ctrl_inst.latch_mem_inst.RAM\[24\]\[6\]
+ sky130_fd_sc_hd__and3_2
XFILLER_0_16_166 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[28\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[28\]\[5\] net202 dig_ctrl_inst.latch_mem_inst.gclk\[28\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[17\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[17\]\[3\] net217 dig_ctrl_inst.latch_mem_inst.gclk\[17\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_77_309 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
Xhold90 VGND VDPWR VDPWR VGND net372 net22 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_169 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1576_ VDPWR VGND VDPWR VGND _0285_ _0286_ _0284_ _0288_ sky130_fd_sc_hd__or3_4
X_1645_ VDPWR VGND VDPWR VGND _0356_ net72 net121 dig_ctrl_inst.latch_mem_inst.RAM\[14\]\[1\]
+ sky130_fd_sc_hd__and3_2
X_1714_ VDPWR VGND VDPWR VGND _0135_ dig_ctrl_inst.latch_mem_inst.RAM\[31\]\[2\] _0132_
+ _0424_ dig_ctrl_inst.latch_mem_inst.RAM\[33\]\[2\] sky130_fd_sc_hd__a22o_1
Xrebuffer11 VDPWR VGND VDPWR VGND net293 _1028_ sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_0_67_52 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xrebuffer22 VDPWR VGND VDPWR VGND net304 _1076_ sky130_fd_sc_hd__buf_2
X_2128_ VGND VDPWR VDPWR VGND _0820_ net171 _0819_ net168 _0813_ sky130_fd_sc_hd__a211o_1
X_2059_ VDPWR VGND VDPWR VGND _0752_ _0751_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_180 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_42_209 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[28\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[28\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[28\] sky130_fd_sc_hd__clkbuf_4
X_1430_ VDPWR VGND VDPWR VGND net254 dig_ctrl_inst.cpu_inst.r0\[7\] net259 _0171_
+ sky130_fd_sc_hd__or3_1
X_1292_ VGND VDPWR VDPWR VGND net136 _1136_ net135 sky130_fd_sc_hd__and2_4
X_1361_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[36\] net57 net97
+ net154 sky130_fd_sc_hd__and3_2
XFILLER_0_68_3 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_1628_ VGND VDPWR VDPWR VGND _0339_ net52 net99 net102 dig_ctrl_inst.latch_mem_inst.RAM\[39\]\[1\]
+ sky130_fd_sc_hd__and4_1
X_1559_ VGND VDPWR VDPWR VGND _0272_ _0237_ _0269_ _0271_ net252 _0270_ sky130_fd_sc_hd__o2111ai_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[61\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[61\]\[5\] net199 dig_ctrl_inst.latch_mem_inst.gclk\[61\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_61_Left_139 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[50\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[50\]\[3\] net215 dig_ctrl_inst.latch_mem_inst.gclk\[50\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_70_Left_148 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_32_253 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_23_57 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xrebuffer2 VDPWR VGND VDPWR VGND net284 net283 sky130_fd_sc_hd__dlygate4sd1_1
X_2393_ VGND VDPWR VDPWR VGND clknet_leaf_4_clk net341 net179 dig_ctrl_inst.synchronizer_port_i_inst\[0\].out
+ sky130_fd_sc_hd__dfrtp_1
X_2462_ VGND VDPWR VDPWR VGND clknet_leaf_3_clk net335 net173 dig_ctrl_inst.mode_sync
+ sky130_fd_sc_hd__dfrtp_1
X_1413_ VDPWR VGND VDPWR VGND dig_ctrl_inst.cpu_inst.rst_ni _0161_ sky130_fd_sc_hd__inv_2
X_2531_ VDPWR VGND VDPWR VGND uio_out[4] net277 sky130_fd_sc_hd__buf_2
XFILLER_0_2_125 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1275_ VGND VDPWR VDPWR VGND net267 _1123_ dig_ctrl_inst.cpu_inst.r2\[4\] sky130_fd_sc_hd__and2b_1
X_1344_ VDPWR VGND VDPWR VGND _0130_ net69 _1140_ net106 sky130_fd_sc_hd__and3_2
XFILLER_0_61_337 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xfanout177 VGND VDPWR VDPWR VGND net180 net177 sky130_fd_sc_hd__clkbuf_4
Xfanout133 VGND VDPWR VDPWR VGND _1063_ net133 sky130_fd_sc_hd__clkbuf_4
Xfanout144 VGND VDPWR VDPWR VGND net147 net144 sky130_fd_sc_hd__clkbuf_2
Xfanout166 VDPWR VGND VDPWR VGND net166 _1060_ sky130_fd_sc_hd__buf_2
Xfanout188 VDPWR VGND VDPWR VGND net188 net189 sky130_fd_sc_hd__buf_2
Xfanout155 VGND VDPWR VDPWR VGND net156 net155 sky130_fd_sc_hd__clkbuf_2
Xfanout111 VDPWR VGND VDPWR VGND net111 net112 sky130_fd_sc_hd__buf_2
Xfanout122 VDPWR VGND VDPWR VGND net122 _1128_ sky130_fd_sc_hd__buf_2
Xfanout100 VDPWR VGND VDPWR VGND _1136_ net100 sky130_fd_sc_hd__buf_4
Xfanout199 VGND VDPWR VDPWR VGND net200 net199 sky130_fd_sc_hd__clkbuf_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[54\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[54\]\[4\] net211 dig_ctrl_inst.latch_mem_inst.gclk\[54\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_29_Right_29 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_38_Right_38 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[43\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[43\]\[2\] net227 dig_ctrl_inst.latch_mem_inst.gclk\[43\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_47_Right_47 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[32\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[32\]\[0\] net243 dig_ctrl_inst.latch_mem_inst.gclk\[32\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_56_Right_56 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1962_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[27\]\[6\] _0130_ _0668_
+ _0142_ dig_ctrl_inst.latch_mem_inst.RAM\[42\]\[6\] _0663_ sky130_fd_sc_hd__a221o_1
XFILLER_0_43_337 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1893_ VDPWR VGND VDPWR VGND _0129_ dig_ctrl_inst.latch_mem_inst.RAM\[2\]\[5\] _1133_
+ _0600_ dig_ctrl_inst.latch_mem_inst.RAM\[26\]\[5\] sky130_fd_sc_hd__a22o_1
XFILLER_0_11_212 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_2514_ VGND VDPWR VDPWR VGND clknet_leaf_9_clk _0111_ net141 dig_ctrl_inst.cpu_inst.cpu_state\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_2376_ VGND VDPWR VDPWR VGND clknet_leaf_4_clk _0003_ net177 dig_ctrl_inst.spi_receiver_inst.spi_cnt\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_65_Right_65 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_59_97 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_2445_ VGND VDPWR VDPWR VGND clknet_leaf_11_clk _0053_ net140 dig_ctrl_inst.cpu_inst.r1\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_1258_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.r1\[5\] net263 _1106_ net267
+ sky130_fd_sc_hd__and3b_1
X_1189_ VDPWR VGND VDPWR VGND _1037_ net170 sky130_fd_sc_hd__inv_2
X_1327_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[18\] net61 net109
+ net148 sky130_fd_sc_hd__and3_2
XPHY_EDGE_ROW_74_Right_74 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[20\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[20\]\[7\] net185 dig_ctrl_inst.latch_mem_inst.gclk\[20\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_46_120 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_61_178 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[58\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[58\]\[5\] net205 dig_ctrl_inst.latch_mem_inst.gclk\[58\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[47\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[47\]\[3\] net220 dig_ctrl_inst.latch_mem_inst.gclk\[47\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[36\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[36\]\[1\] net236 dig_ctrl_inst.latch_mem_inst.gclk\[36\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_29_23 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
X_2230_ VGND VDPWR VDPWR VGND _0747_ _0918_ _0912_ sky130_fd_sc_hd__nand2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[2\].gen_latches\[7\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[2\]\[7\] net186 dig_ctrl_inst.latch_mem_inst.gclk\[2\]
+ sky130_fd_sc_hd__dlxtp_1
X_2092_ VDPWR VGND VDPWR VGND _0785_ _1014_ _0745_ sky130_fd_sc_hd__or2_2
X_2161_ VGND VDPWR VDPWR VGND _0255_ _0258_ _0254_ _0852_ sky130_fd_sc_hd__o21a_1
XFILLER_0_43_101 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_28_131 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_1945_ VGND VDPWR VDPWR VGND _0651_ net65 net91 net117 dig_ctrl_inst.latch_mem_inst.RAM\[25\]\[6\]
+ sky130_fd_sc_hd__and4_1
XFILLER_0_43_156 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_1876_ VGND VDPWR VDPWR VGND _0583_ net62 net103 net131 dig_ctrl_inst.latch_mem_inst.RAM\[19\]\[5\]
+ sky130_fd_sc_hd__and4_1
X_2359_ VGND VDPWR VDPWR VGND _0108_ net372 _0988_ dig_ctrl_inst.cpu_inst.port_o\[5\]
+ sky130_fd_sc_hd__mux2_1
X_2428_ VGND VDPWR VDPWR VGND clknet_leaf_9_clk _0036_ net142 dig_ctrl_inst.cpu_inst.data\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[13\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[13\]\[6\] net192 dig_ctrl_inst.latch_mem_inst.gclk\[13\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_8_Left_86 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_31_46 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1730_ VGND VDPWR VDPWR VGND _0440_ net70 net79 dig_ctrl_inst.latch_mem_inst.RAM\[28\]\[2\]
+ _0120_ dig_ctrl_inst.latch_mem_inst.RAM\[17\]\[2\] sky130_fd_sc_hd__a32o_1
XFILLER_0_40_104 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1592_ VDPWR VGND VDPWR VGND _0304_ _1138_ net122 dig_ctrl_inst.latch_mem_inst.RAM\[6\]\[0\]
+ sky130_fd_sc_hd__and3_2
XFILLER_0_31_79 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1661_ VGND VDPWR VDPWR VGND _0372_ net44 net103 net131 dig_ctrl_inst.latch_mem_inst.RAM\[51\]\[1\]
+ sky130_fd_sc_hd__and4_1
X_2144_ VGND VDPWR VDPWR VGND _0046_ _0835_ net41 dig_ctrl_inst.cpu_inst.r0\[1\] sky130_fd_sc_hd__mux2_1
X_2213_ VGND VDPWR VDPWR VGND _0902_ _1125_ _0878_ sky130_fd_sc_hd__or2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[29\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[29\]\[0\] net243 dig_ctrl_inst.latch_mem_inst.gclk\[29\]
+ sky130_fd_sc_hd__dlxtp_1
X_2075_ VDPWR VGND VDPWR VGND _0742_ _0744_ net163 _0768_ sky130_fd_sc_hd__or3_4
X_1928_ VDPWR VGND VDPWR VGND _0634_ net65 net77 dig_ctrl_inst.latch_mem_inst.RAM\[28\]\[6\]
+ sky130_fd_sc_hd__and3_2
X_1859_ VGND VDPWR VDPWR VGND _0030_ _0565_ _0276_ net253 sky130_fd_sc_hd__mux2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[17\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[17\]\[7\] net187 dig_ctrl_inst.latch_mem_inst.gclk\[17\]
+ sky130_fd_sc_hd__dlxtp_1
Xhold91 VGND VDPWR VDPWR VGND net373 dig_ctrl_inst.cpu_inst.r3\[2\] sky130_fd_sc_hd__dlygate4sd3_1
Xhold80 VGND VDPWR VDPWR VGND net362 dig_ctrl_inst.cpu_inst.r2\[1\] sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_9_109 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1713_ VDPWR VGND VDPWR VGND _0420_ _0422_ _0421_ _0404_ _0423_ sky130_fd_sc_hd__or4_1
XFILLER_0_5_337 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1575_ VGND VDPWR VDPWR VGND _0286_ _0284_ _0287_ _0285_ sky130_fd_sc_hd__nor3_4
X_1644_ VDPWR VGND VDPWR VGND _0355_ net109 net120 dig_ctrl_inst.latch_mem_inst.RAM\[2\]\[1\]
+ sky130_fd_sc_hd__and3_2
Xrebuffer23 VGND VDPWR VDPWR VGND net305 net304 sky130_fd_sc_hd__clkbuf_1
X_2127_ VDPWR VGND VDPWR VGND _0819_ _0818_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_3 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2058_ VGND VDPWR VDPWR VGND _0751_ _0746_ _0749_ _0747_ _0743_ sky130_fd_sc_hd__or4b_4
X_1360_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[35\] net148 _0137_
+ sky130_fd_sc_hd__and2_1
X_1291_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[3\] net155 _1135_
+ sky130_fd_sc_hd__and2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[62\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[62\]\[0\] net244 dig_ctrl_inst.latch_mem_inst.gclk\[62\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[10\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[10\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[10\] clknet_leaf_0_clk sky130_fd_sc_hd__dlclkp_1
X_1627_ VGND VDPWR VDPWR VGND _0026_ _0338_ _0276_ net268 sky130_fd_sc_hd__mux2_1
X_1558_ VGND VDPWR VDPWR VGND _0233_ _0172_ _0271_ sky130_fd_sc_hd__nand2b_1
X_1489_ VGND VDPWR VDPWR VGND _0207_ dig_ctrl_inst.cpu_inst.data\[1\] _0198_ net161
+ sky130_fd_sc_hd__mux2_1
X_2519__269 VGND VDPWR VDPWR VGND net269 _2519__269/HI sky130_fd_sc_hd__conb_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[50\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[50\]\[7\] net183 dig_ctrl_inst.latch_mem_inst.gclk\[50\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_2_3 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_2530_ VDPWR VGND VDPWR VGND uio_out[3] net276 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_21_Left_99 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xrebuffer3 VDPWR VGND VDPWR VGND net285 net283 sky130_fd_sc_hd__dlygate4sd1_1
X_2392_ VGND VDPWR VDPWR VGND clknet_leaf_4_clk net3 net175 dig_ctrl_inst.synchronizer_port_i_inst\[0\].pipe\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_2461_ VGND VDPWR VDPWR VGND clknet_leaf_3_clk net14 net173 dig_ctrl_inst.synchronizer_mode_i_inst.pipe\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_1412_ VGND VDPWR VDPWR VGND _0161_ _1002_ net180 sky130_fd_sc_hd__nand2_2
X_1343_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[26\] net70 net83
+ net153 sky130_fd_sc_hd__and3_2
X_1274_ VDPWR VGND VDPWR VGND _1122_ dig_ctrl_inst.cpu_inst.r3\[4\] net264 net267
+ sky130_fd_sc_hd__and3_2
Xwire36 VGND VDPWR VDPWR VGND net36 _0621_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_16_clk VGND VDPWR VDPWR VGND clknet_leaf_16_clk clknet_1_0__leaf_clk
+ sky130_fd_sc_hd__clkbuf_8
Xfanout178 VDPWR VGND VDPWR VGND net178 net180 sky130_fd_sc_hd__buf_2
Xfanout101 VGND VDPWR VDPWR VGND _1136_ net101 sky130_fd_sc_hd__clkbuf_4
Xfanout123 VDPWR VGND VDPWR VGND net123 net127 sky130_fd_sc_hd__buf_2
Xfanout145 VGND VDPWR VDPWR VGND net146 net145 sky130_fd_sc_hd__clkbuf_4
Xfanout189 VDPWR VGND VDPWR VGND net189 net190 sky130_fd_sc_hd__buf_2
Xfanout156 VGND VDPWR VDPWR VGND _1097_ net156 sky130_fd_sc_hd__clkbuf_2
Xfanout112 VGND VDPWR VDPWR VGND net113 net112 sky130_fd_sc_hd__clkbuf_2
Xfanout167 VDPWR VGND VDPWR VGND net167 net168 sky130_fd_sc_hd__buf_2
XFILLER_0_64_176 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[43\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[43\]\[6\] net193 dig_ctrl_inst.latch_mem_inst.gclk\[43\]
+ sky130_fd_sc_hd__dlxtp_1
X_1892_ VDPWR VGND VDPWR VGND _0157_ dig_ctrl_inst.latch_mem_inst.RAM\[24\]\[5\] _0127_
+ _0599_ dig_ctrl_inst.latch_mem_inst.RAM\[60\]\[5\] sky130_fd_sc_hd__a22o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[32\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[32\]\[4\] net211 dig_ctrl_inst.latch_mem_inst.gclk\[32\]
+ sky130_fd_sc_hd__dlxtp_1
X_1961_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[9\]\[6\] _1143_ _0667_
+ _0148_ dig_ctrl_inst.latch_mem_inst.RAM\[49\]\[6\] _0660_ sky130_fd_sc_hd__a221o_1
X_2513_ VGND VDPWR VDPWR VGND clknet_leaf_5_clk _0110_ net179 net24 sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_5_clk VGND VDPWR VDPWR VGND clknet_leaf_5_clk clknet_1_1__leaf_clk sky130_fd_sc_hd__clkbuf_8
X_2375_ VGND VDPWR VDPWR VGND clknet_leaf_5_clk _0002_ net177 dig_ctrl_inst.spi_receiver_inst.spi_cnt\[0\]
+ sky130_fd_sc_hd__dfrtp_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[21\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[21\]\[2\] net226 dig_ctrl_inst.latch_mem_inst.gclk\[21\]
+ sky130_fd_sc_hd__dlxtp_1
X_1326_ VDPWR VGND VDPWR VGND _0121_ net111 net65 sky130_fd_sc_hd__and2_1
X_2444_ VGND VDPWR VDPWR VGND clknet_leaf_11_clk _0052_ net142 dig_ctrl_inst.cpu_inst.r0\[7\]
+ sky130_fd_sc_hd__dfrtp_2
X_1257_ VGND VDPWR VDPWR VGND _1105_ _1010_ _1025_ _1103_ sky130_fd_sc_hd__and3_4
X_1188_ VGND VDPWR VDPWR VGND _1018_ _1032_ _1033_ _1034_ _1035_ _1036_ sky130_fd_sc_hd__o41a_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[59\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[59\]\[0\] net244 dig_ctrl_inst.latch_mem_inst.gclk\[59\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_46_165 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[10\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[10\]\[0\] net240 dig_ctrl_inst.latch_mem_inst.gclk\[10\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_37_132 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[47\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[47\]\[7\] net189 dig_ctrl_inst.latch_mem_inst.gclk\[47\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[3\].gen_latches\[2\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[3\]\[2\] net231 dig_ctrl_inst.latch_mem_inst.gclk\[3\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_29_57 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2160_ VDPWR VGND VDPWR VGND _0851_ _0850_ _0848_ _0845_ sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[36\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[36\]\[5\] net206 dig_ctrl_inst.latch_mem_inst.gclk\[36\]
+ sky130_fd_sc_hd__dlxtp_1
X_2091_ VGND VDPWR VDPWR VGND net161 _0784_ _0783_ sky130_fd_sc_hd__nand2_1
X_1875_ VGND VDPWR VDPWR VGND _1139_ dig_ctrl_inst.latch_mem_inst.RAM\[7\]\[5\] _0579_
+ _0580_ _0581_ _0582_ sky130_fd_sc_hd__a2111o_1
X_1944_ VGND VDPWR VDPWR VGND _0650_ net45 net81 net104 dig_ctrl_inst.latch_mem_inst.RAM\[63\]\[6\]
+ sky130_fd_sc_hd__and4_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[25\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[25\]\[3\] net216 dig_ctrl_inst.latch_mem_inst.gclk\[25\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_9_12 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2427_ VGND VDPWR VDPWR VGND clknet_leaf_9_clk _0035_ net141 dig_ctrl_inst.cpu_inst.data\[1\]
+ sky130_fd_sc_hd__dfrtp_2
Xdig_ctrl_inst.latch_mem_inst.gen_input_latches\[3\].n_latch VGND VDPWR VDPWR VGND
+ dig_ctrl_inst.latch_mem_inst.wdata\[3\] dig_ctrl_inst.data_out\[3\] clknet_leaf_8_clk
+ sky130_fd_sc_hd__dlxtn_1
X_2358_ VGND VDPWR VDPWR VGND _0107_ net21 _0988_ dig_ctrl_inst.cpu_inst.port_o\[4\]
+ sky130_fd_sc_hd__mux2_1
X_2289_ VGND VDPWR VDPWR VGND _0880_ _0877_ _0971_ _0751_ sky130_fd_sc_hd__o21ai_1
X_1309_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[11\] net155 _1145_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_43_3 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
Xdig_ctrl_inst.latch_mem_inst.gen_words\[14\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[14\]\[1\] net235 dig_ctrl_inst.latch_mem_inst.gclk\[14\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_74_293 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[7\].gen_latches\[3\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[7\]\[3\] net222 dig_ctrl_inst.latch_mem_inst.gclk\[7\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[15\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[15\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[15\] clknet_leaf_1_clk sky130_fd_sc_hd__dlclkp_1
X_1660_ VGND VDPWR VDPWR VGND _0371_ net101 net108 net127 dig_ctrl_inst.latch_mem_inst.RAM\[7\]\[1\]
+ sky130_fd_sc_hd__and4_1
X_1591_ VDPWR VGND VDPWR VGND _0303_ net45 net94 dig_ctrl_inst.latch_mem_inst.RAM\[54\]\[0\]
+ sky130_fd_sc_hd__and3_2
X_2212_ VGND VDPWR VDPWR VGND _1125_ _0901_ _0878_ sky130_fd_sc_hd__nand2_1
X_2143_ VDPWR VGND VDPWR VGND _0753_ _0830_ _0835_ _0834_ _0755_ _0833_ sky130_fd_sc_hd__a221o_1
XFILLER_0_56_77 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_72_32 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[29\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[29\]\[4\] net214 dig_ctrl_inst.latch_mem_inst.gclk\[29\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_8_324 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2074_ VGND VDPWR VDPWR VGND _1068_ _0760_ _0264_ _0766_ _0767_ sky130_fd_sc_hd__o22a_1
XFILLER_0_12_330 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_1858_ VDPWR VGND VDPWR VGND _0566_ _0565_ sky130_fd_sc_hd__inv_2
X_1927_ VGND VDPWR VDPWR VGND _0633_ net55 net99 net103 dig_ctrl_inst.latch_mem_inst.RAM\[39\]\[6\]
+ sky130_fd_sc_hd__and4_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[31\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[31\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[31\] sky130_fd_sc_hd__clkbuf_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[18\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[18\]\[2\] net226 dig_ctrl_inst.latch_mem_inst.gclk\[18\]
+ sky130_fd_sc_hd__dlxtp_1
X_1789_ VGND VDPWR VDPWR VGND _0114_ dig_ctrl_inst.latch_mem_inst.RAM\[13\]\[3\] _0495_
+ _0496_ _0497_ _0498_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_26_25 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xhold70 VGND VDPWR VDPWR VGND net352 dig_ctrl_inst.cpu_inst.r3\[6\] sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 VGND VDPWR VDPWR VGND net363 dig_ctrl_inst.cpu_inst.r2\[6\] sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 VGND VDPWR VDPWR VGND net374 dig_ctrl_inst.cpu_inst.r1\[0\] sky130_fd_sc_hd__dlygate4sd3_1
X_1712_ VDPWR VGND VDPWR VGND _0278_ dig_ctrl_inst.latch_mem_inst.RAM\[9\]\[2\] _1143_
+ _0422_ dig_ctrl_inst.latch_mem_inst.RAM\[5\]\[2\] sky130_fd_sc_hd__a22o_1
XANTENNA_1 VGND VDPWR VDPWR VGND _0325_ sky130_fd_sc_hd__diode_2
X_1643_ VDPWR VGND VDPWR VGND _0354_ net63 net87 dig_ctrl_inst.latch_mem_inst.RAM\[24\]\[1\]
+ sky130_fd_sc_hd__and3_2
X_1574_ VDPWR VGND VDPWR VGND _0117_ _0116_ _1148_ _1143_ _0286_ sky130_fd_sc_hd__or4_4
X_2126_ VGND VDPWR VDPWR VGND _0768_ _0816_ _0817_ _0765_ _0818_ sky130_fd_sc_hd__o22ai_1
X_2057_ VDPWR VGND VDPWR VGND _0750_ _1011_ net283 sky130_fd_sc_hd__or2_2
Xrebuffer13 VDPWR VGND VDPWR VGND net295 _1073_ sky130_fd_sc_hd__dlygate4sd1_1
X_1290_ VGND VDPWR VDPWR VGND _1135_ net132 net126 net106 sky130_fd_sc_hd__and3_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[62\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[62\]\[4\] net214 dig_ctrl_inst.latch_mem_inst.gclk\[62\]
+ sky130_fd_sc_hd__dlxtp_1
X_1626_ VDPWR VGND VDPWR VGND _0338_ _0324_ _0326_ _0337_ dig_ctrl_inst.latch_mem_inst.RAM\[0\]\[0\]
+ _0288_ sky130_fd_sc_hd__o32a_1
XFILLER_0_5_113 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[51\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[51\]\[2\] net229 dig_ctrl_inst.latch_mem_inst.gclk\[51\]
+ sky130_fd_sc_hd__dlxtp_1
X_1557_ VGND VDPWR VDPWR VGND _0270_ _0236_ _0167_ net138 sky130_fd_sc_hd__nand3b_1
X_1488_ VGND VDPWR VDPWR VGND _0019_ dig_ctrl_inst.cpu_inst.ip\[0\] _0204_ _0206_
+ sky130_fd_sc_hd__mux2_1
X_2109_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.data\[0\] _0802_ _0800_ _0801_
+ sky130_fd_sc_hd__and3b_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[40\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[40\]\[0\] net244 dig_ctrl_inst.latch_mem_inst.gclk\[40\]
+ sky130_fd_sc_hd__dlxtp_1
X_2460_ VGND VDPWR VDPWR VGND clknet_leaf_11_clk _0068_ net140 dig_ctrl_inst.cpu_inst.r2\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xrebuffer4 VDPWR VGND VDPWR VGND net286 net283 sky130_fd_sc_hd__dlygate4sd1_1
X_2391_ VGND VDPWR VDPWR VGND clknet_leaf_4_clk net342 net179 dig_ctrl_inst.synchronizer_port_i_inst\[1\].out
+ sky130_fd_sc_hd__dfrtp_1
X_1273_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.r1\[4\] net263 _1121_ net267
+ sky130_fd_sc_hd__and3b_1
X_1342_ VDPWR VGND VDPWR VGND net83 net69 _0129_ sky130_fd_sc_hd__and2_2
X_1411_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[63\] net152 _0160_
+ sky130_fd_sc_hd__and2_1
Xwire37 VGND VDPWR VDPWR VGND net37 net38 sky130_fd_sc_hd__clkbuf_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[24\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[24\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[24\] sky130_fd_sc_hd__clkbuf_4
X_1609_ VGND VDPWR VDPWR VGND _0321_ net58 net72 dig_ctrl_inst.latch_mem_inst.RAM\[46\]\[0\]
+ _0138_ dig_ctrl_inst.latch_mem_inst.RAM\[37\]\[0\] sky130_fd_sc_hd__a32o_1
Xfanout102 VDPWR VGND VDPWR VGND net105 net102 sky130_fd_sc_hd__buf_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[55\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[55\]\[3\] net216 dig_ctrl_inst.latch_mem_inst.gclk\[55\]
+ sky130_fd_sc_hd__dlxtp_1
Xfanout179 VGND VDPWR VDPWR VGND net180 net179 sky130_fd_sc_hd__clkbuf_4
Xfanout135 VDPWR VGND VDPWR VGND _1062_ net135 sky130_fd_sc_hd__buf_4
Xfanout146 VDPWR VGND VDPWR VGND net146 net147 sky130_fd_sc_hd__buf_2
Xfanout124 VGND VDPWR VDPWR VGND net125 net124 sky130_fd_sc_hd__clkbuf_2
Xfanout168 VDPWR VGND VDPWR VGND net168 _1054_ sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout157 VDPWR VGND VDPWR VGND net157 net158 sky130_fd_sc_hd__buf_2
X_2532__278 VGND VDPWR VDPWR VGND net278 _2532__278/HI sky130_fd_sc_hd__conb_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[44\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[44\]\[1\] net234 dig_ctrl_inst.latch_mem_inst.gclk\[44\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_20_247 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1960_ VDPWR VGND VDPWR VGND _0644_ _0648_ _0646_ _0656_ _0666_ sky130_fd_sc_hd__or4_4
X_1891_ VDPWR VGND VDPWR VGND _0595_ _0597_ _0596_ _0594_ _0598_ sky130_fd_sc_hd__or4_1
X_2512_ VGND VDPWR VDPWR VGND clknet_leaf_5_clk _0109_ net179 net23 sky130_fd_sc_hd__dfrtp_1
X_2443_ VGND VDPWR VDPWR VGND clknet_leaf_10_clk _0051_ net142 dig_ctrl_inst.cpu_inst.r0\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[22\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[22\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[22\] clknet_leaf_17_clk sky130_fd_sc_hd__dlclkp_1
X_2374_ VDPWR VGND VDPWR VGND net282 net2 dig_ctrl_inst.latch_mem_inst.rst_ni sky130_fd_sc_hd__dfxtp_1
X_1325_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[17\] net155 _0120_
+ sky130_fd_sc_hd__and2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[21\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[21\]\[6\] net198 dig_ctrl_inst.latch_mem_inst.gclk\[21\]
+ sky130_fd_sc_hd__dlxtp_1
X_1256_ VDPWR VGND VDPWR VGND _1104_ _1103_ sky130_fd_sc_hd__inv_2
X_1187_ VDPWR VGND VDPWR VGND net256 dig_ctrl_inst.cpu_inst.r0\[3\] net260 _1035_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_61_169 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_61_136 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[59\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[59\]\[4\] net214 dig_ctrl_inst.latch_mem_inst.gclk\[59\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_49_Left_127 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_46_155 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[10\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[10\]\[4\] net208 dig_ctrl_inst.latch_mem_inst.gclk\[10\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_6_285 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_339 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_58_Left_136 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[48\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[48\]\[2\] net225 dig_ctrl_inst.latch_mem_inst.gclk\[48\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_67_Left_145 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_76_Left_154 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[3\].gen_latches\[6\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[3\]\[6\] net196 dig_ctrl_inst.latch_mem_inst.gclk\[3\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[37\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[37\]\[0\] net245 dig_ctrl_inst.latch_mem_inst.gclk\[37\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_52_136 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_20_49 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_46 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_2090_ VGND VDPWR VDPWR VGND net254 net258 _1015_ _0783_ sky130_fd_sc_hd__nor3b_4
XFILLER_0_0_15 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_1943_ VDPWR VGND VDPWR VGND _0649_ net88 net125 dig_ctrl_inst.latch_mem_inst.RAM\[8\]\[6\]
+ sky130_fd_sc_hd__and3_2
X_1874_ VDPWR VGND VDPWR VGND _0581_ net59 net97 dig_ctrl_inst.latch_mem_inst.RAM\[36\]\[5\]
+ sky130_fd_sc_hd__and3_2
XFILLER_0_28_155 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_2426_ VGND VDPWR VDPWR VGND clknet_leaf_8_clk _0034_ net143 dig_ctrl_inst.cpu_inst.data\[0\]
+ sky130_fd_sc_hd__dfrtp_4
Xdig_ctrl_inst.latch_mem_inst.gen_input_latches\[7\].n_latch VGND VDPWR VDPWR VGND
+ dig_ctrl_inst.latch_mem_inst.wdata\[7\] dig_ctrl_inst.data_out\[7\] clknet_leaf_8_clk
+ sky130_fd_sc_hd__dlxtn_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[25\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[25\]\[7\] net189 dig_ctrl_inst.latch_mem_inst.gclk\[25\]
+ sky130_fd_sc_hd__dlxtp_1
X_2357_ VGND VDPWR VDPWR VGND _0106_ net386 _0988_ dig_ctrl_inst.cpu_inst.port_o\[3\]
+ sky130_fd_sc_hd__mux2_1
X_1308_ VGND VDPWR VDPWR VGND _1145_ net106 net126 net92 sky130_fd_sc_hd__and3_4
X_2288_ VGND VDPWR VDPWR VGND _0055_ _0970_ _0967_ net369 sky130_fd_sc_hd__mux2_1
X_1239_ VDPWR VGND VDPWR VGND _1087_ dig_ctrl_inst.cpu_inst.r3\[1\] net262 net266
+ sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[14\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[14\]\[5\] net201 dig_ctrl_inst.latch_mem_inst.gclk\[14\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[7\].gen_latches\[7\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[7\]\[7\] net188 dig_ctrl_inst.latch_mem_inst.gclk\[7\]
+ sky130_fd_sc_hd__dlxtp_1
X_1590_ VDPWR VGND VDPWR VGND _0302_ net48 net78 dig_ctrl_inst.latch_mem_inst.RAM\[60\]\[0\]
+ sky130_fd_sc_hd__and3_2
XFILLER_0_56_23 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_0_225 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_2142_ VDPWR VGND VDPWR VGND _0804_ dig_ctrl_inst.synchronizer_port_i_inst\[1\].out
+ _0802_ _0834_ dig_ctrl_inst.spi_data_o\[1\] sky130_fd_sc_hd__a22o_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[17\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[17\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[17\] sky130_fd_sc_hd__clkbuf_4
X_2211_ VGND VDPWR VDPWR VGND _0900_ _0788_ _0885_ _0889_ _0899_ sky130_fd_sc_hd__o211a_1
X_2073_ VGND VDPWR VDPWR VGND net161 _0766_ _0759_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_336 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
X_1857_ VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[0\]\[4\] _0288_ _0564_
+ _0519_ _0565_ sky130_fd_sc_hd__o22a_2
XFILLER_0_12_320 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1788_ VDPWR VGND VDPWR VGND _0497_ net87 net122 dig_ctrl_inst.latch_mem_inst.RAM\[8\]\[3\]
+ sky130_fd_sc_hd__and3_2
X_1926_ VGND VDPWR VDPWR VGND _0632_ net43 net80 net116 dig_ctrl_inst.latch_mem_inst.RAM\[61\]\[6\]
+ sky130_fd_sc_hd__and4_1
X_2409_ VGND VDPWR VDPWR VGND clknet_leaf_5_clk _0017_ net145 dig_ctrl_inst.cpu_inst.port_o\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[18\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[18\]\[6\] net197 dig_ctrl_inst.latch_mem_inst.gclk\[18\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_22_128 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_180 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xhold60 VGND VDPWR VDPWR VGND net342 dig_ctrl_inst.synchronizer_port_i_inst\[1\].pipe\[0\]
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 VGND VDPWR VDPWR VGND net353 net24 sky130_fd_sc_hd__dlygate4sd3_1
Xhold93 VGND VDPWR VDPWR VGND net375 dig_ctrl_inst.cpu_inst.r1\[3\] sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 VGND VDPWR VDPWR VGND net364 dig_ctrl_inst.cpu_inst.r3\[7\] sky130_fd_sc_hd__dlygate4sd3_1
X_1711_ VGND VDPWR VDPWR VGND _0421_ net70 net74 dig_ctrl_inst.latch_mem_inst.RAM\[30\]\[2\]
+ _0142_ dig_ctrl_inst.latch_mem_inst.RAM\[42\]\[2\] sky130_fd_sc_hd__a32o_1
XANTENNA_2 VGND VDPWR VDPWR VGND _0443_ sky130_fd_sc_hd__diode_2
X_1642_ VDPWR VGND VDPWR VGND _0353_ net64 net96 dig_ctrl_inst.latch_mem_inst.RAM\[20\]\[1\]
+ sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[1\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[1\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[1\] clknet_leaf_19_clk sky130_fd_sc_hd__dlclkp_1
X_1573_ VGND VDPWR VDPWR VGND net119 net132 _1133_ _1142_ _0277_ _0285_ sky130_fd_sc_hd__a2111o_1
X_2125_ VGND VDPWR VDPWR VGND _0817_ net157 _0779_ sky130_fd_sc_hd__or2_1
X_2056_ VGND VDPWR VDPWR VGND _1011_ net284 _0749_ sky130_fd_sc_hd__nor2_1
Xrebuffer14 VDPWR VGND VDPWR VGND net296 dig_ctrl_inst.cpu_inst.instr\[4\] sky130_fd_sc_hd__dlygate4sd1_1
X_1909_ VDPWR VGND VDPWR VGND _0616_ net61 net128 dig_ctrl_inst.latch_mem_inst.RAM\[16\]\[5\]
+ sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[27\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[27\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[27\] clknet_leaf_1_clk sky130_fd_sc_hd__dlclkp_1
XFILLER_0_53_57 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_5_136 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1625_ VDPWR VGND VDPWR VGND _0320_ _0336_ _0331_ _0287_ _0337_ sky130_fd_sc_hd__or4_1
X_1556_ VDPWR VGND VDPWR VGND _0269_ _1119_ net159 _0244_ _1104_ net160 sky130_fd_sc_hd__o32a_1
X_1487_ VGND VDPWR VDPWR VGND _0206_ _0205_ _0173_ _1001_ sky130_fd_sc_hd__mux2_1
X_2039_ VGND VDPWR VDPWR VGND _0035_ _0398_ _0741_ dig_ctrl_inst.cpu_inst.data\[1\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_109 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_30_Left_108 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[51\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[51\]\[6\] net192 dig_ctrl_inst.latch_mem_inst.gclk\[51\]
+ sky130_fd_sc_hd__dlxtp_1
X_2108_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.data\[2\] _0801_ dig_ctrl_inst.cpu_inst.data\[3\]
+ sky130_fd_sc_hd__nor2_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[40\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[40\]\[4\] net208 dig_ctrl_inst.latch_mem_inst.gclk\[40\]
+ sky130_fd_sc_hd__dlxtp_1
X_1410_ VDPWR VGND VDPWR VGND _0160_ net50 net82 net108 sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[63\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[63\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[63\] sky130_fd_sc_hd__clkbuf_4
Xrebuffer5 VDPWR VGND VDPWR VGND net287 net286 sky130_fd_sc_hd__dlymetal6s2s_1
X_2390_ VGND VDPWR VDPWR VGND clknet_leaf_4_clk net4 net175 dig_ctrl_inst.synchronizer_port_i_inst\[1\].pipe\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_1272_ VDPWR VGND VDPWR VGND _1120_ _1118_ _1025_ _1010_ sky130_fd_sc_hd__and3_2
XFILLER_0_64_45 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
X_1341_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[25\] net148 _0128_
+ sky130_fd_sc_hd__and2_1
Xwire38 VGND VDPWR VDPWR VGND net38 _0578_ sky130_fd_sc_hd__clkbuf_1
Xfanout147 VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.rst_ni net147 sky130_fd_sc_hd__clkbuf_2
Xfanout125 VGND VDPWR VDPWR VGND net127 net125 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_66_3 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_1608_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[8\]\[0\] _1142_ _0320_
+ _0153_ dig_ctrl_inst.latch_mem_inst.RAM\[55\]\[0\] _0319_ sky130_fd_sc_hd__a221o_1
X_1539_ VGND VDPWR VDPWR VGND _0249_ _0252_ _0251_ sky130_fd_sc_hd__nand2_1
Xfanout103 VGND VDPWR VDPWR VGND net105 net103 sky130_fd_sc_hd__clkbuf_2
Xfanout114 VDPWR VGND VDPWR VGND net115 net114 sky130_fd_sc_hd__buf_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[55\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[55\]\[7\] net184 dig_ctrl_inst.latch_mem_inst.gclk\[55\]
+ sky130_fd_sc_hd__dlxtp_1
Xfanout169 VDPWR VGND VDPWR VGND net169 _1045_ sky130_fd_sc_hd__buf_2
Xfanout158 VDPWR VGND VDPWR VGND net158 _1067_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_49_175 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
Xdig_ctrl_inst.latch_mem_inst.gen_words\[0\].gen_latches\[0\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[0\]\[0\] net246 dig_ctrl_inst.latch_mem_inst.gclk\[0\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[44\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[44\]\[5\] net200 dig_ctrl_inst.latch_mem_inst.gclk\[44\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_37_337 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[33\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[33\]\[3\] net215 dig_ctrl_inst.latch_mem_inst.gclk\[33\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_16_Right_16 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_55_134 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
Xdig_ctrl_inst.latch_mem_inst.gen_words\[22\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[22\]\[1\] net236 dig_ctrl_inst.latch_mem_inst.gclk\[22\]
+ sky130_fd_sc_hd__dlxtp_1
X_1890_ VGND VDPWR VDPWR VGND _0597_ net64 net77 dig_ctrl_inst.latch_mem_inst.RAM\[28\]\[5\]
+ _0154_ dig_ctrl_inst.latch_mem_inst.RAM\[57\]\[5\] sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_25_Right_25 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2511_ VGND VDPWR VDPWR VGND clknet_leaf_5_clk _0108_ net179 net22 sky130_fd_sc_hd__dfrtp_1
X_2442_ VGND VDPWR VDPWR VGND clknet_leaf_6_clk _0050_ net145 dig_ctrl_inst.cpu_inst.r0\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_2373_ VGND VDPWR VDPWR VGND _0990_ _0996_ _0201_ _0113_ sky130_fd_sc_hd__o21a_1
X_1186_ VGND VDPWR VDPWR VGND net260 _1034_ dig_ctrl_inst.cpu_inst.r2\[3\] sky130_fd_sc_hd__and2b_1
X_1255_ VGND VDPWR VDPWR VGND _1103_ _1102_ _1101_ _1100_ _1099_ _1018_ sky130_fd_sc_hd__o41a_4
X_1324_ VGND VDPWR VDPWR VGND _0120_ net132 net119 net71 sky130_fd_sc_hd__and3_4
XPHY_EDGE_ROW_34_Right_34 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_19_337 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_43_Right_43 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_6_297 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_6_253 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_52_Right_52 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[4\].gen_latches\[1\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[4\]\[1\] net237 dig_ctrl_inst.latch_mem_inst.gclk\[4\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[48\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[48\]\[6\] net192 dig_ctrl_inst.latch_mem_inst.gclk\[48\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_61_Right_61 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_52_148 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_37_189 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_70_Right_70 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[37\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[37\]\[4\] net208 dig_ctrl_inst.latch_mem_inst.gclk\[37\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[6\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[6\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[6\] clknet_leaf_17_clk sky130_fd_sc_hd__dlclkp_1
X_1942_ VGND VDPWR VDPWR VGND _0648_ net107 net124 net132 dig_ctrl_inst.latch_mem_inst.RAM\[3\]\[6\]
+ sky130_fd_sc_hd__and4_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[26\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[26\]\[2\] net230 dig_ctrl_inst.latch_mem_inst.gclk\[26\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_61_57 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
X_1873_ VGND VDPWR VDPWR VGND _0580_ net59 net101 net107 dig_ctrl_inst.latch_mem_inst.RAM\[39\]\[5\]
+ sky130_fd_sc_hd__and4_1
XFILLER_0_28_178 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2356_ VGND VDPWR VDPWR VGND _0105_ net385 _0988_ dig_ctrl_inst.cpu_inst.port_o\[2\]
+ sky130_fd_sc_hd__mux2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[15\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[15\]\[0\] net243 dig_ctrl_inst.latch_mem_inst.gclk\[15\]
+ sky130_fd_sc_hd__dlxtp_1
X_2425_ VGND VDPWR VDPWR VGND clknet_leaf_13_clk _0033_ net139 dig_ctrl_inst.cpu_inst.instr\[7\]
+ sky130_fd_sc_hd__dfrtp_2
X_2287_ VGND VDPWR VDPWR VGND _0856_ _0854_ _0970_ _0751_ sky130_fd_sc_hd__o21ai_1
X_1307_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[10\] net83 net124
+ net154 sky130_fd_sc_hd__and3_2
XFILLER_0_29_3 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_1238_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.r1\[1\] net262 _1086_ net266
+ sky130_fd_sc_hd__and3b_1
X_1169_ VDPWR VGND VDPWR VGND net252 dig_ctrl_inst.cpu_inst.instr\[6\] net253 dig_ctrl_inst.cpu_inst.instr\[7\]
+ _1017_ sky130_fd_sc_hd__or4_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[8\].gen_latches\[2\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[8\]\[2\] net225 dig_ctrl_inst.latch_mem_inst.gclk\[8\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[56\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[56\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[56\] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_237 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_2210_ VGND VDPWR VDPWR VGND _0899_ _0750_ _0892_ _0893_ _0898_ sky130_fd_sc_hd__o211a_1
XFILLER_0_0_204 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_12 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_2072_ VGND VDPWR VDPWR VGND _0765_ net163 _0764_ sky130_fd_sc_hd__nand2_2
X_2141_ VGND VDPWR VDPWR VGND _0820_ _0822_ _0833_ _0832_ sky130_fd_sc_hd__nand3_1
X_1925_ VDPWR VGND VDPWR VGND _0631_ net43 net110 dig_ctrl_inst.latch_mem_inst.RAM\[50\]\[6\]
+ sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[34\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[34\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[34\] clknet_leaf_17_clk sky130_fd_sc_hd__dlclkp_1
X_1856_ VDPWR VGND VDPWR VGND _0563_ _0558_ _0551_ _0534_ _0564_ sky130_fd_sc_hd__or4_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[19\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[19\]\[1\] net239 dig_ctrl_inst.latch_mem_inst.gclk\[19\]
+ sky130_fd_sc_hd__dlxtp_1
X_1787_ VGND VDPWR VDPWR VGND _0496_ net56 net91 net104 dig_ctrl_inst.latch_mem_inst.RAM\[43\]\[3\]
+ sky130_fd_sc_hd__and4_1
X_2408_ VGND VDPWR VDPWR VGND clknet_leaf_6_clk _0016_ net145 dig_ctrl_inst.cpu_inst.port_o\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_2339_ VGND VDPWR VDPWR VGND _0090_ dig_ctrl_inst.spi_data_i\[3\] _0986_ dig_ctrl_inst.cpu_inst.port_o\[3\]
+ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_2_Right_2 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_62_232 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xhold61 VGND VDPWR VDPWR VGND net343 dig_ctrl_inst.stb_d sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 VGND VDPWR VDPWR VGND net354 dig_ctrl_inst.cpu_inst.prev_state\[2\] sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 VGND VDPWR VDPWR VGND net376 dig_ctrl_inst.cpu_inst.r3\[4\] sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 VGND VDPWR VDPWR VGND net365 dig_ctrl_inst.cpu_inst.r1\[5\] sky130_fd_sc_hd__dlygate4sd3_1
Xhold50 VGND VDPWR VDPWR VGND net332 dig_ctrl_inst.synchronizer_port_i_inst\[4\].pipe\[0\]
+ sky130_fd_sc_hd__dlygate4sd3_1
X_1572_ VDPWR VGND VDPWR VGND _0281_ _0283_ _0282_ _0280_ _0284_ sky130_fd_sc_hd__or4_2
XANTENNA_3 VGND VDPWR VDPWR VGND _0477_ sky130_fd_sc_hd__diode_2
X_1710_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[21\]\[2\] _0124_ _0420_
+ _0151_ dig_ctrl_inst.latch_mem_inst.RAM\[53\]\[2\] _0415_ sky130_fd_sc_hd__a221o_1
X_1641_ VGND VDPWR VDPWR VGND _0352_ net62 net99 net116 dig_ctrl_inst.latch_mem_inst.RAM\[21\]\[1\]
+ sky130_fd_sc_hd__and4_1
XFILLER_0_6_48 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2124_ VGND VDPWR VDPWR VGND _0814_ _0815_ _0816_ sky130_fd_sc_hd__nor2_1
Xrebuffer15 VDPWR VGND VDPWR VGND _1026_ net297 sky130_fd_sc_hd__buf_6
X_2055_ VGND VDPWR VDPWR VGND _0748_ _1015_ _1031_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_101 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1839_ VDPWR VGND VDPWR VGND _0547_ net58 net111 dig_ctrl_inst.latch_mem_inst.RAM\[34\]\[4\]
+ sky130_fd_sc_hd__and3_2
XFILLER_0_32_70 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
X_1908_ VGND VDPWR VDPWR VGND _0158_ dig_ctrl_inst.latch_mem_inst.RAM\[61\]\[5\] _0612_
+ _0613_ _0614_ _0615_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_12_29 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[63\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[63\]\[3\] net220 dig_ctrl_inst.latch_mem_inst.gclk\[63\]
+ sky130_fd_sc_hd__dlxtp_1
X_1624_ VDPWR VGND VDPWR VGND _0333_ _0335_ _0334_ _0332_ _0336_ sky130_fd_sc_hd__or4_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[52\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[52\]\[1\] net239 dig_ctrl_inst.latch_mem_inst.gclk\[52\]
+ sky130_fd_sc_hd__dlxtp_1
X_1555_ VGND VDPWR VDPWR VGND _0245_ _0267_ _0268_ sky130_fd_sc_hd__nor2_1
X_2107_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.data\[1\] _0799_ _0800_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_19_clk VGND VDPWR VDPWR VGND clknet_leaf_19_clk clknet_1_1__leaf_clk
+ sky130_fd_sc_hd__clkbuf_8
X_1486_ VGND VDPWR VDPWR VGND _0205_ dig_ctrl_inst.cpu_inst.data\[0\] _0198_ net164
+ sky130_fd_sc_hd__mux2_1
X_2038_ VGND VDPWR VDPWR VGND _0034_ _0338_ _0741_ dig_ctrl_inst.cpu_inst.data\[0\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_313 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_17_221 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_4_192 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[49\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[49\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[49\] sky130_fd_sc_hd__clkbuf_4
Xrebuffer6 VDPWR VGND VDPWR VGND net288 net287 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_0_48_25 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1340_ VDPWR VGND VDPWR VGND _0128_ net61 net90 net114 sky130_fd_sc_hd__and3_2
X_1271_ VDPWR VGND VDPWR VGND _1119_ _1118_ sky130_fd_sc_hd__inv_2
Xwire39 VGND VDPWR VDPWR VGND net39 net40 sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_8_clk VGND VDPWR VDPWR VGND clknet_leaf_8_clk clknet_1_1__leaf_clk sky130_fd_sc_hd__clkbuf_8
Xdig_ctrl_inst.latch_mem_inst.gen_words\[56\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[56\]\[2\] net229 dig_ctrl_inst.latch_mem_inst.gclk\[56\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_38_80 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xfanout126 VGND VDPWR VDPWR VGND net127 net126 sky130_fd_sc_hd__clkbuf_2
X_1469_ VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_addr\[5\] _0186_ _0195_ _0197_ sky130_fd_sc_hd__or3b_1
Xfanout148 VGND VDPWR VDPWR VGND net151 net148 sky130_fd_sc_hd__clkbuf_2
X_1538_ VGND VDPWR VDPWR VGND _0251_ net170 net169 sky130_fd_sc_hd__or2_1
X_1607_ VDPWR VGND VDPWR VGND _0150_ dig_ctrl_inst.latch_mem_inst.RAM\[51\]\[0\] _0149_
+ _0319_ dig_ctrl_inst.latch_mem_inst.RAM\[52\]\[0\] sky130_fd_sc_hd__a22o_1
Xfanout104 VDPWR VGND VDPWR VGND net104 net105 sky130_fd_sc_hd__buf_2
Xfanout159 VDPWR VGND VDPWR VGND net159 _1125_ sky130_fd_sc_hd__buf_2
Xfanout115 VDPWR VGND VDPWR VGND net116 net115 sky130_fd_sc_hd__buf_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[45\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[45\]\[0\] net243 dig_ctrl_inst.latch_mem_inst.gclk\[45\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[0\].gen_latches\[4\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[0\]\[4\] net211 dig_ctrl_inst.latch_mem_inst.gclk\[0\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_0_3 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_113 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[33\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[33\]\[7\] net183 dig_ctrl_inst.latch_mem_inst.gclk\[33\]
+ sky130_fd_sc_hd__dlxtp_1
X_2510_ VGND VDPWR VDPWR VGND clknet_leaf_5_clk _0107_ net179 net21 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_48 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_50_59 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[39\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[39\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[39\] clknet_leaf_2_clk sky130_fd_sc_hd__dlclkp_1
X_2441_ VGND VDPWR VDPWR VGND clknet_leaf_6_clk _0049_ net145 dig_ctrl_inst.cpu_inst.r0\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[22\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[22\]\[5\] net200 dig_ctrl_inst.latch_mem_inst.gclk\[22\]
+ sky130_fd_sc_hd__dlxtp_1
X_2372_ VGND VDPWR VDPWR VGND _0112_ dig_ctrl_inst.cpu_inst.cpu_state\[1\] _0990_
+ _1027_ sky130_fd_sc_hd__mux2_1
X_1323_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[16\] net62 net150
+ net128 sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[11\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[11\]\[3\] net222 dig_ctrl_inst.latch_mem_inst.gclk\[11\]
+ sky130_fd_sc_hd__dlxtp_1
X_1185_ VGND VDPWR VDPWR VGND net257 _1033_ dig_ctrl_inst.cpu_inst.r1\[3\] sky130_fd_sc_hd__and2b_1
X_1254_ VDPWR VGND VDPWR VGND net257 dig_ctrl_inst.cpu_inst.r0\[5\] net260 _1102_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_6_243 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[49\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[49\]\[1\] net237 dig_ctrl_inst.latch_mem_inst.gclk\[49\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_6_265 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[20\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[20\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[20\] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_260 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[41\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[41\]._gclk
+ dig_ctrl_inst.latch_mem_inst.data_we\[41\] clknet_leaf_13_clk sky130_fd_sc_hd__dlclkp_1
XFILLER_0_4_81 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[6\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[6\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[6\] sky130_fd_sc_hd__clkbuf_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[4\].gen_latches\[5\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[4\]\[5\] net204 dig_ctrl_inst.latch_mem_inst.gclk\[4\]
+ sky130_fd_sc_hd__dlxtp_1
X_1941_ VGND VDPWR VDPWR VGND _0647_ net48 net92 net107 dig_ctrl_inst.latch_mem_inst.RAM\[59\]\[6\]
+ sky130_fd_sc_hd__and4_1
X_1872_ VDPWR VGND VDPWR VGND _0579_ net59 net83 dig_ctrl_inst.latch_mem_inst.RAM\[42\]\[5\]
+ sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[26\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[26\]\[6\] net194 dig_ctrl_inst.latch_mem_inst.gclk\[26\]
+ sky130_fd_sc_hd__dlxtp_1
X_2355_ VGND VDPWR VDPWR VGND _0104_ net392 _0988_ dig_ctrl_inst.cpu_inst.port_o\[1\]
+ sky130_fd_sc_hd__mux2_1
X_1306_ VGND VDPWR VDPWR VGND net290 _1144_ net136 _1062_ _1078_ net134 sky130_fd_sc_hd__a2111oi_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[15\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[15\]\[4\] net214 dig_ctrl_inst.latch_mem_inst.gclk\[15\]
+ sky130_fd_sc_hd__dlxtp_1
X_2424_ VGND VDPWR VDPWR VGND clknet_leaf_13_clk _0032_ net139 dig_ctrl_inst.cpu_inst.instr\[6\]
+ sky130_fd_sc_hd__dfrtp_2
X_2286_ VGND VDPWR VDPWR VGND _0054_ _0969_ _0967_ net367 sky130_fd_sc_hd__mux2_1
X_1237_ VDPWR VGND VDPWR VGND _1085_ net163 _1025_ _1010_ sky130_fd_sc_hd__and3_2
XFILLER_0_19_113 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1168_ VGND VDPWR VDPWR VGND _1016_ net252 net253 sky130_fd_sc_hd__or2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[8\].gen_latches\[6\].p_latch VGND VDPWR VDPWR
+ VGND dig_ctrl_inst.latch_mem_inst.RAM\[8\]\[6\] net196 dig_ctrl_inst.latch_mem_inst.gclk\[8\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_0_216 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_2140_ VDPWR VGND VDPWR VGND _0832_ _0831_ _0827_ _0824_ _0787_ _0257_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_0_249 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_72_24 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2071_ VGND VDPWR VDPWR VGND _0742_ _0744_ _0764_ sky130_fd_sc_hd__nor2_1
X_1855_ VDPWR VGND VDPWR VGND _0560_ _0562_ _0561_ _0559_ _0563_ sky130_fd_sc_hd__or4_1
X_1924_ VDPWR VGND VDPWR VGND _0630_ net50 net84 dig_ctrl_inst.latch_mem_inst.RAM\[58\]\[6\]
+ sky130_fd_sc_hd__and3_2
XFILLER_0_16_116 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1786_ VGND VDPWR VDPWR VGND _0495_ net71 net82 net119 dig_ctrl_inst.latch_mem_inst.RAM\[29\]\[3\]
+ sky130_fd_sc_hd__and4_1
XFILLER_0_12_300 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
Xdig_ctrl_inst.latch_mem_inst.gen_words\[19\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[19\]\[5\] net200 dig_ctrl_inst.latch_mem_inst.gclk\[19\]
+ sky130_fd_sc_hd__dlxtp_1
X_2338_ VGND VDPWR VDPWR VGND _0089_ dig_ctrl_inst.spi_data_i\[2\] _0986_ dig_ctrl_inst.cpu_inst.port_o\[2\]
+ sky130_fd_sc_hd__mux2_1
X_2407_ VGND VDPWR VDPWR VGND clknet_leaf_6_clk _0015_ net145 dig_ctrl_inst.cpu_inst.port_o\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_3 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
X_2269_ VGND VDPWR VDPWR VGND _0955_ net170 _0860_ net167 _0954_ sky130_fd_sc_hd__a211o_1
XFILLER_0_39_208 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_1_82 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xhold40 VGND VDPWR VDPWR VGND net322 dig_ctrl_inst.latch_mem_inst.wdata\[6\] sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 VGND VDPWR VDPWR VGND net333 dig_ctrl_inst.spi_receiver_inst.synchronizer_spi_sclk.pipe\[0\]
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 VGND VDPWR VDPWR VGND net355 dig_ctrl_inst.spi_miso_o sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 VGND VDPWR VDPWR VGND net366 dig_ctrl_inst.cpu_inst.r2\[5\] sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 VGND VDPWR VDPWR VGND net344 dig_ctrl_inst.spi_receiver_inst.spi_sclk_sync
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_16 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
Xhold95 VGND VDPWR VDPWR VGND net377 dig_ctrl_inst.cpu_inst.r1\[7\] sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_49 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
X_1571_ VDPWR VGND VDPWR VGND _0283_ net92 net123 _1093_ sky130_fd_sc_hd__and3_2
X_1640_ VGND VDPWR VDPWR VGND _0351_ net56 net81 net104 dig_ctrl_inst.latch_mem_inst.RAM\[47\]\[1\]
+ sky130_fd_sc_hd__and4_1
XANTENNA_4 VGND VDPWR VDPWR VGND _0511_ sky130_fd_sc_hd__diode_2
X_2123_ VGND VDPWR VDPWR VGND net157 _0775_ _0815_ sky130_fd_sc_hd__nor2_1
Xrebuffer16 VDPWR VGND VDPWR VGND net298 net181 sky130_fd_sc_hd__dlymetal6s2s_1
X_2054_ VGND VDPWR VDPWR VGND _1031_ _0747_ _1015_ sky130_fd_sc_hd__nor2_2
X_1838_ VGND VDPWR VDPWR VGND _0139_ dig_ctrl_inst.latch_mem_inst.RAM\[39\]\[4\] _0543_
+ _0544_ _0545_ _0546_ sky130_fd_sc_hd__a2111o_1
Xdig_ctrl_inst.latch_mem_inst.gen_gclk\[13\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gen_gclk\[13\]._gclk
+ dig_ctrl_inst.latch_mem_inst.gclk\[13\] sky130_fd_sc_hd__clkbuf_4
X_1907_ VDPWR VGND VDPWR VGND _0614_ net76 net120 dig_ctrl_inst.latch_mem_inst.RAM\[12\]\[5\]
+ sky130_fd_sc_hd__and3_2
X_1769_ VDPWR VGND VDPWR VGND _0478_ net44 net128 dig_ctrl_inst.latch_mem_inst.RAM\[48\]\[3\]
+ sky130_fd_sc_hd__and3_2
Xoutput30 VDPWR VGND VDPWR VGND uo_out[2] net30 sky130_fd_sc_hd__buf_2
XFILLER_0_35_277 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_37_16 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[63\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[63\]\[7\] net185 dig_ctrl_inst.latch_mem_inst.gclk\[63\]
+ sky130_fd_sc_hd__dlxtp_1
X_1623_ VGND VDPWR VDPWR VGND _1139_ dig_ctrl_inst.latch_mem_inst.RAM\[7\]\[0\] _0290_
+ _0300_ _0301_ _0335_ sky130_fd_sc_hd__a2111o_1
X_1554_ VGND VDPWR VDPWR VGND _0253_ _0265_ net169 _1037_ _0267_ _0266_ sky130_fd_sc_hd__o221a_1
X_1485_ VGND VDPWR VDPWR VGND _0204_ _0201_ _0203_ _0199_ _1030_ sky130_fd_sc_hd__or4b_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[52\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[52\]\[5\] net201 dig_ctrl_inst.latch_mem_inst.gclk\[52\]
+ sky130_fd_sc_hd__dlxtp_1
.ends

.subckt res_poly a_n141_4996# a_n141_n5432# VSUBS
X0 a_n141_4996# a_n141_n5432# VSUBS sky130_fd_pr__res_high_po_1p41 l=50.12
.ends

.subckt sky130_leo_ip__rdac_8bit D0 D1 D2 D3 D4 D5 D6 D7 OUT VGND
Xres_poly_0 m1_5556_10930# m1_4470_10930# VGND res_poly
Xres_poly_1 m1_4470_10930# m1_4832_499# VGND res_poly
Xres_poly_2 m1_4470_10930# m1_3384_10930# VGND res_poly
Xres_poly_3 D2 m1_3746_499# VGND res_poly
Xres_poly_4 m1_3384_10930# m1_3746_499# VGND res_poly
Xres_poly_5 m1_3384_10930# m1_2298_10930# VGND res_poly
Xres_poly_6 D1 m1_2660_499# VGND res_poly
Xres_poly_7 m1_2298_10930# m1_2660_499# VGND res_poly
Xres_poly_8 m1_2298_10930# m1_1212_10930# VGND res_poly
Xres_poly_9 VGND m1_1574_499# VGND res_poly
Xres_poly_21 D6 m1_8090_499# VGND res_poly
Xres_poly_20 m1_7728_10930# m1_8090_499# VGND res_poly
Xres_poly_10 m1_1212_10930# m1_1574_499# VGND res_poly
Xres_poly_22 OUT m1_7728_10930# VGND res_poly
Xres_poly_11 m1_1212_10930# m1_850_499# VGND res_poly
Xres_poly_23 OUT m1_9176_499# VGND res_poly
Xres_poly_12 VGND VGND VGND res_poly
Xres_poly_24 D7 m1_9176_499# VGND res_poly
Xres_poly_13 D3 m1_4832_499# VGND res_poly
Xres_poly_25 VGND VGND VGND res_poly
Xres_poly_14 m1_5556_10930# m1_5918_499# VGND res_poly
Xres_poly_15 D4 m1_5918_499# VGND res_poly
Xres_poly_26 D0 m1_850_499# VGND res_poly
Xres_poly_16 m1_6642_10930# m1_5556_10930# VGND res_poly
Xres_poly_18 D5 m1_7004_499# VGND res_poly
Xres_poly_17 m1_6642_10930# m1_7004_499# VGND res_poly
Xres_poly_19 m1_7728_10930# m1_6642_10930# VGND res_poly
.ends

.subckt pfet a_60_n40# w_n242_n247# a_160_0# a_0_0#
X0 a_160_0# a_60_n40# a_0_0# w_n242_n247# sky130_fd_pr__pfet_g5v0d10v5 ad=6 pd=40.6 as=6 ps=40.6 w=20 l=0.5
.ends

.subckt res_poly$1 a_n285_2496# a_n415_n3062# a_n285_n2932#
X0 a_n285_2496# a_n285_n2932# a_n415_n3062# sky130_fd_pr__res_xhigh_po_2p85 l=25.12
.ends

.subckt pfet$10 a_60_n40# w_n242_n247# a_1060_0# a_0_0#
X0 a_1060_0# a_60_n40# a_0_0# w_n242_n247# sky130_fd_pr__pfet_g5v0d10v5 ad=3 pd=20.6 as=3 ps=20.6 w=10 l=5
.ends

.subckt nfet$5 a_60_n40# a_160_0# a_0_0# a_n149_n154#
X0 a_160_0# a_60_n40# a_0_0# a_n149_n154# sky130_fd_pr__nfet_g5v0d10v5 ad=0.3 pd=2.6 as=0.3 ps=2.6 w=1 l=0.5
.ends

.subckt pfet$9 a_60_n40# w_n242_n247# a_1060_0# a_0_0#
X0 a_1060_0# a_60_n40# a_0_0# w_n242_n247# sky130_fd_pr__pfet_g5v0d10v5 ad=0.3 pd=2.6 as=0.3 ps=2.6 w=1 l=5
.ends

.subckt nfet$1 a_60_n40# a_160_0# a_0_0# a_n149_n154#
X0 a_160_0# a_60_n40# a_0_0# a_n149_n154# sky130_fd_pr__nfet_g5v0d10v5 ad=3 pd=20.6 as=3 ps=20.6 w=10 l=0.5
.ends

.subckt sky130_fd_sc_hvl__buf_4$VAR1 VPB VPWR VNB VGND A X
X0 a_149_81# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.21 ps=1.78 w=1.5 l=0.5
X1 VGND a_149_81# X VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X2 X a_149_81# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.21375 ps=2.07 w=0.75 l=0.5
X3 X a_149_81# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X4 VPWR a_149_81# X VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X5 a_149_81# A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.105 ps=1.03 w=0.75 l=0.5
X6 VPWR a_149_81# X VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X7 X a_149_81# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.4275 ps=3.57 w=1.5 l=0.5
X8 X a_149_81# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X9 VGND a_149_81# X VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
.ends

.subckt pfet$5 a_60_n40# w_n242_n247# a_160_0# a_0_0#
X0 a_160_0# a_60_n40# a_0_0# w_n242_n247# sky130_fd_pr__pfet_g5v0d10v5 ad=1.5 pd=10.6 as=1.5 ps=10.6 w=5 l=0.5
.ends

.subckt sky130_fd_sc_hvl__buf_4$1 VPB VPWR VNB VGND A X
X0 a_149_81# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.21 ps=1.78 w=1.5 l=0.5
X1 VGND a_149_81# X VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X2 X a_149_81# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.21375 ps=2.07 w=0.75 l=0.5
X3 X a_149_81# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X4 VPWR a_149_81# X VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X5 a_149_81# A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.105 ps=1.03 w=0.75 l=0.5
X6 VPWR a_149_81# X VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X7 X a_149_81# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.4275 ps=3.57 w=1.5 l=0.5
X8 X a_149_81# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X9 VGND a_149_81# X VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
.ends

.subckt nfet$4 a_60_n40# a_160_0# a_0_0# a_n149_n154#
X0 a_160_0# a_60_n40# a_0_0# a_n149_n154# sky130_fd_pr__nfet_g5v0d10v5 ad=1.5 pd=10.6 as=1.5 ps=10.6 w=5 l=0.5
.ends

.subckt sky130_fd_sc_hvl__nand2_1 VPB VPWR VNB VGND B Y A
X0 a_233_111# B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.07875 pd=0.96 as=0.21375 ps=2.07 w=0.75 l=0.5
X1 Y A a_233_111# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.07875 ps=0.96 w=0.75 l=0.5
X2 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.21 ps=1.78 w=1.5 l=0.5
X3 Y B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.4275 ps=3.57 w=1.5 l=0.5
.ends

.subckt sky130_leo_ip__comparator VDD IN_P OUT_P IN_N CLK OUT_N VSS
Xpfet_0 IN_N VDD m1_1831_3328# m1_1572_726# pfet
Xpfet_1 IN_P VDD COMP_N m1_1831_3328# pfet
Xres_poly$1_0 m1_282_7668# VSS VSS res_poly$1
Xpfet$10_0 m1_282_7668# VDD VDD m1_1831_3328# pfet$10
Xnfet$5_0 COMP_N SR_set VSS VSS nfet$5
Xnfet$5_1 m1_1572_726# SR_reset VSS VSS nfet$5
Xpfet$9_0 m1_282_7668# VDD m1_282_7668# VDD pfet$9
Xnfet$1_0 CLK COMP_N m1_1572_726# VSS nfet$1
Xsky130_fd_sc_hvl__buf_4$VAR1_0 VDD VDD VSS VSS sky130_fd_sc_hvl__nand2_1_1/Y OUT_N
+ sky130_fd_sc_hvl__buf_4$VAR1
Xpfet$5_0 COMP_N VDD VDD SR_set pfet$5
Xpfet$5_1 m1_1572_726# VDD VDD SR_reset pfet$5
Xsky130_fd_sc_hvl__buf_4$1_0 VDD VDD VSS VSS sky130_fd_sc_hvl__nand2_1_1/A OUT_P sky130_fd_sc_hvl__buf_4$1
Xnfet$4_0 COMP_N m1_1572_726# VSS VSS nfet$4
Xsky130_fd_sc_hvl__nand2_1_0 VDD VDD VSS VSS sky130_fd_sc_hvl__nand2_1_1/Y sky130_fd_sc_hvl__nand2_1_1/A
+ SR_reset sky130_fd_sc_hvl__nand2_1
Xnfet$4_1 m1_1572_726# VSS COMP_N VSS nfet$4
Xsky130_fd_sc_hvl__nand2_1_1 VDD VDD VSS VSS SR_set sky130_fd_sc_hvl__nand2_1_1/Y
+ sky130_fd_sc_hvl__nand2_1_1/A sky130_fd_sc_hvl__nand2_1
.ends

.subckt tt_um_tt08_aicd_playground VAPWR ui_in[7] ui_in[6] ui_in[5] ui_in[4] ui_in[3]
+ ui_in[2] ui_in[1] ui_in[0] VDPWR VGND uio_in[7] uio_in[6] uio_in[5] uio_in[4] uio_in[3]
+ uio_in[2] uio_in[1] uio_in[0] ena uo_out[7] uo_out[6] uo_out[5] uo_out[4] uo_out[3]
+ uo_out[2] uo_out[1] uo_out[0] clk rst_n uio_out[7] uio_out[6] uio_out[5] uio_out[4]
+ uio_out[3] uio_out[2] uio_out[1] uio_out[0] uio_oe[7] uio_oe[6] uio_oe[5] uio_oe[4]
+ uio_oe[3] uio_oe[2] uio_oe[1] uio_oe[0] ua[7] ua[6] ua[5] ua[4] ua[3] ua[2] ua[1]
+ ua[0]
Xsky130_leo_ip__levelshifter_up_1 VAPWR VDPWR sky130_fd_sc_hvl__buf_4_1/A dig_ctrl_top_0/port_ms_o[6]
+ VGND sky130_leo_ip__levelshifter_up
Xsky130_leo_ip__levelshifter_up_2 VAPWR VDPWR sky130_fd_sc_hvl__buf_4_2/A dig_ctrl_top_0/port_ms_o[5]
+ VGND sky130_leo_ip__levelshifter_up
Xsky130_leo_ip__levelshifter_up_3 VAPWR VDPWR sky130_fd_sc_hvl__buf_4_3/A dig_ctrl_top_0/port_ms_o[4]
+ VGND sky130_leo_ip__levelshifter_up
Xsky130_leo_ip__levelshifter_up_4 VAPWR VDPWR sky130_fd_sc_hvl__buf_4_4/A dig_ctrl_top_0/port_ms_o[3]
+ VGND sky130_leo_ip__levelshifter_up
Xsky130_leo_ip__levelshifter_up_5 VAPWR VDPWR sky130_fd_sc_hvl__buf_4_5/A dig_ctrl_top_0/port_ms_o[2]
+ VGND sky130_leo_ip__levelshifter_up
Xsky130_fd_sc_hvl__buf_4_0 VGND VGND VAPWR VAPWR sky130_fd_sc_hvl__buf_4_0/X sky130_fd_sc_hvl__buf_4_0/A
+ sky130_fd_sc_hvl__buf_4
Xsky130_leo_ip__levelshifter_up_6 VAPWR VDPWR sky130_fd_sc_hvl__buf_4_6/A dig_ctrl_top_0/port_ms_o[1]
+ VGND sky130_leo_ip__levelshifter_up
Xsky130_fd_sc_hvl__buf_4_1 VGND VGND VAPWR VAPWR sky130_fd_sc_hvl__buf_4_1/X sky130_fd_sc_hvl__buf_4_1/A
+ sky130_fd_sc_hvl__buf_4
Xsky130_leo_ip__levelshifter_up_7 VAPWR VDPWR sky130_fd_sc_hvl__buf_4_7/A dig_ctrl_top_0/port_ms_o[0]
+ VGND sky130_leo_ip__levelshifter_up
Xsky130_fd_sc_hvl__buf_4_2 VGND VGND VAPWR VAPWR sky130_fd_sc_hvl__buf_4_2/X sky130_fd_sc_hvl__buf_4_2/A
+ sky130_fd_sc_hvl__buf_4
Xsky130_leo_ip__levelshifter_down_0 VDPWR dig_ctrl_top_0/port_ms_i sky130_leo_ip__comparator_0/OUT_P
+ VGND sky130_leo_ip__levelshifter_down
Xdig_ctrl_top_0 uio_in[4] clk ena rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4]
+ ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[5] uio_in[6]
+ uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6]
+ uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6]
+ uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6]
+ uo_out[7] dig_ctrl_top_0/clk_o dig_ctrl_top_0/port_ms_i dig_ctrl_top_0/port_ms_o[0]
+ dig_ctrl_top_0/port_ms_o[1] dig_ctrl_top_0/port_ms_o[2] dig_ctrl_top_0/port_ms_o[3]
+ dig_ctrl_top_0/port_ms_o[4] dig_ctrl_top_0/port_ms_o[5] dig_ctrl_top_0/port_ms_o[6]
+ dig_ctrl_top_0/port_ms_o[7] VDPWR VGND dig_ctrl_top
Xsky130_fd_sc_hvl__buf_4_4 VGND VGND VAPWR VAPWR sky130_fd_sc_hvl__buf_4_4/X sky130_fd_sc_hvl__buf_4_4/A
+ sky130_fd_sc_hvl__buf_4
Xsky130_fd_sc_hvl__buf_4_3 VGND VGND VAPWR VAPWR sky130_fd_sc_hvl__buf_4_3/X sky130_fd_sc_hvl__buf_4_3/A
+ sky130_fd_sc_hvl__buf_4
Xsky130_fd_sc_hvl__buf_4_5 VGND VGND VAPWR VAPWR sky130_fd_sc_hvl__buf_4_5/X sky130_fd_sc_hvl__buf_4_5/A
+ sky130_fd_sc_hvl__buf_4
Xsky130_fd_sc_hvl__buf_4_6 VGND VGND VAPWR VAPWR sky130_fd_sc_hvl__buf_4_6/X sky130_fd_sc_hvl__buf_4_6/A
+ sky130_fd_sc_hvl__buf_4
Xsky130_fd_sc_hvl__buf_4_7 VGND VGND VAPWR VAPWR sky130_fd_sc_hvl__buf_4_7/X sky130_fd_sc_hvl__buf_4_7/A
+ sky130_fd_sc_hvl__buf_4
Xsky130_leo_ip__rdac_8bit_0 sky130_fd_sc_hvl__buf_4_7/X sky130_fd_sc_hvl__buf_4_6/X
+ sky130_fd_sc_hvl__buf_4_5/X sky130_fd_sc_hvl__buf_4_4/X sky130_fd_sc_hvl__buf_4_3/X
+ sky130_fd_sc_hvl__buf_4_2/X sky130_fd_sc_hvl__buf_4_1/X sky130_fd_sc_hvl__buf_4_0/X
+ ua[1] VGND sky130_leo_ip__rdac_8bit
Xsky130_leo_ip__comparator_0 VAPWR ua[0] sky130_leo_ip__comparator_0/OUT_P ua[1] dig_ctrl_top_0/clk_o
+ sky130_leo_ip__comparator_0/OUT_N VGND sky130_leo_ip__comparator
Xsky130_leo_ip__levelshifter_up_0 VAPWR VDPWR sky130_fd_sc_hvl__buf_4_0/A dig_ctrl_top_0/port_ms_o[7]
+ VGND sky130_leo_ip__levelshifter_up
.ends

