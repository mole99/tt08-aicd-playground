VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_tt08_aicd_playground
  CLASS BLOCK ;
  FOREIGN tt_um_tt08_aicd_playground ;
  ORIGIN 0.000 0.000 ;
  SIZE 319.240 BY 225.760 ;
  PIN VDPWR
    ANTENNADIFFAREA 6.800000 ;
    PORT
      LAYER met4 ;
        RECT 181.200 6.240 182.800 221.625 ;
    END
    PORT
      LAYER met4 ;
        RECT 197.400 6.240 199.000 218.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 21.040 6.240 22.640 218.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 141.040 6.240 142.640 218.880 ;
    END
  END VDPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 184.000 6.240 185.600 221.625 ;
    END
    PORT
      LAYER met4 ;
        RECT 200.200 6.240 201.800 218.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 24.340 6.240 25.940 218.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 144.340 6.240 145.940 218.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 312.200 6.240 313.800 218.880 ;
    END
  END VGND
  PIN VAPWR
    ANTENNADIFFAREA 4.016000 ;
    PORT
      LAYER met4 ;
        RECT 190.000 6.240 191.600 221.625 ;
    END
    PORT
      LAYER met4 ;
        RECT 203.000 6.240 204.600 218.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 315.000 6.240 316.600 218.880 ;
    END
  END VAPWR
  PIN clk
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met4 ;
        RECT 128.190 224.760 128.490 225.760 ;
    END
  END clk
  PIN ena
    PORT
      LAYER met4 ;
        RECT 130.950 224.760 131.250 225.760 ;
    END
  END ena
  PIN rst_n
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END rst_n
  PIN ua[0]
    ANTENNAGATEAREA 0.710000 ;
    ANTENNADIFFAREA 1.260000 ;
    PORT
      LAYER met4 ;
        RECT 136.170 0.000 137.070 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    ANTENNAGATEAREA 10.000000 ;
    PORT
      LAYER met4 ;
        RECT 116.850 0.000 117.750 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    PORT
      LAYER met4 ;
        RECT 97.530 0.000 98.430 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    PORT
      LAYER met4 ;
        RECT 78.210 0.000 79.110 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    PORT
      LAYER met4 ;
        RECT 58.890 0.000 59.790 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    PORT
      LAYER met4 ;
        RECT 39.570 0.000 40.470 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    PORT
      LAYER met4 ;
        RECT 20.250 0.000 21.150 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    PORT
      LAYER met4 ;
        RECT 0.930 0.000 1.830 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 122.670 224.760 122.970 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 119.910 224.760 120.210 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 117.150 224.760 117.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 111.630 224.760 111.930 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 108.870 224.760 109.170 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 106.110 224.760 106.410 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 100.590 224.760 100.890 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 97.830 224.760 98.130 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    PORT
      LAYER met4 ;
        RECT 95.070 224.760 95.370 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 89.550 224.760 89.850 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    PORT
      LAYER met4 ;
        RECT 86.790 224.760 87.090 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    PORT
      LAYER met4 ;
        RECT 84.030 224.760 84.330 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 34.350 224.760 34.650 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 31.590 224.760 31.890 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 28.830 224.760 29.130 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 23.310 224.760 23.610 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 20.550 224.760 20.850 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 17.790 224.760 18.090 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 56.430 224.760 56.730 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 53.670 224.760 53.970 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 50.910 224.760 51.210 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 45.390 224.760 45.690 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 42.630 224.760 42.930 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 39.870 224.760 40.170 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 78.510 224.760 78.810 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 75.750 224.760 76.050 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 72.990 224.760 73.290 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 67.470 224.760 67.770 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 64.710 224.760 65.010 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 61.950 224.760 62.250 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uo_out[7]
  OBS
      LAYER li1 ;
        RECT 5.520 6.395 313.800 222.085 ;
      LAYER met1 ;
        RECT 1.910 5.840 313.800 223.020 ;
      LAYER met2 ;
        RECT 1.930 0.715 313.800 223.050 ;
      LAYER met3 ;
        RECT 1.905 0.715 317.025 221.625 ;
      LAYER met4 ;
        RECT 3.055 224.360 14.630 224.760 ;
        RECT 15.730 224.360 17.390 224.760 ;
        RECT 18.490 224.360 20.150 224.760 ;
        RECT 21.250 224.360 22.910 224.760 ;
        RECT 24.010 224.360 25.670 224.760 ;
        RECT 26.770 224.360 28.430 224.760 ;
        RECT 29.530 224.360 31.190 224.760 ;
        RECT 32.290 224.360 33.950 224.760 ;
        RECT 35.050 224.360 36.710 224.760 ;
        RECT 37.810 224.360 39.470 224.760 ;
        RECT 40.570 224.360 42.230 224.760 ;
        RECT 43.330 224.360 44.990 224.760 ;
        RECT 46.090 224.360 47.750 224.760 ;
        RECT 48.850 224.360 50.510 224.760 ;
        RECT 51.610 224.360 53.270 224.760 ;
        RECT 54.370 224.360 56.030 224.760 ;
        RECT 57.130 224.360 58.790 224.760 ;
        RECT 59.890 224.360 61.550 224.760 ;
        RECT 62.650 224.360 64.310 224.760 ;
        RECT 65.410 224.360 67.070 224.760 ;
        RECT 68.170 224.360 69.830 224.760 ;
        RECT 70.930 224.360 72.590 224.760 ;
        RECT 73.690 224.360 75.350 224.760 ;
        RECT 76.450 224.360 78.110 224.760 ;
        RECT 79.210 224.360 80.870 224.760 ;
        RECT 81.970 224.360 83.630 224.760 ;
        RECT 84.730 224.360 86.390 224.760 ;
        RECT 87.490 224.360 89.150 224.760 ;
        RECT 90.250 224.360 91.910 224.760 ;
        RECT 93.010 224.360 94.670 224.760 ;
        RECT 95.770 224.360 97.430 224.760 ;
        RECT 98.530 224.360 100.190 224.760 ;
        RECT 101.290 224.360 102.950 224.760 ;
        RECT 104.050 224.360 105.710 224.760 ;
        RECT 106.810 224.360 108.470 224.760 ;
        RECT 109.570 224.360 111.230 224.760 ;
        RECT 112.330 224.360 113.990 224.760 ;
        RECT 115.090 224.360 116.750 224.760 ;
        RECT 117.850 224.360 119.510 224.760 ;
        RECT 120.610 224.360 122.270 224.760 ;
        RECT 123.370 224.360 125.030 224.760 ;
        RECT 126.130 224.360 127.790 224.760 ;
        RECT 128.890 224.360 130.550 224.760 ;
        RECT 131.650 224.360 317.025 224.760 ;
        RECT 3.055 222.025 317.025 224.360 ;
        RECT 3.055 219.280 180.800 222.025 ;
        RECT 3.055 5.840 20.640 219.280 ;
        RECT 23.040 5.840 23.940 219.280 ;
        RECT 26.340 5.840 140.640 219.280 ;
        RECT 143.040 5.840 143.940 219.280 ;
        RECT 146.340 5.840 180.800 219.280 ;
        RECT 183.200 5.840 183.600 222.025 ;
        RECT 186.000 5.840 189.600 222.025 ;
        RECT 192.000 219.280 317.025 222.025 ;
        RECT 192.000 5.840 197.000 219.280 ;
        RECT 199.400 5.840 199.800 219.280 ;
        RECT 202.200 5.840 202.600 219.280 ;
        RECT 205.000 5.840 311.800 219.280 ;
        RECT 314.200 5.840 314.600 219.280 ;
        RECT 317.000 5.840 317.025 219.280 ;
        RECT 3.055 1.400 317.025 5.840 ;
        RECT 3.055 0.715 19.850 1.400 ;
        RECT 21.550 0.715 39.170 1.400 ;
        RECT 40.870 0.715 58.490 1.400 ;
        RECT 60.190 0.715 77.810 1.400 ;
        RECT 79.510 0.715 97.130 1.400 ;
        RECT 98.830 0.715 116.450 1.400 ;
        RECT 118.150 0.715 135.770 1.400 ;
        RECT 137.470 0.715 317.025 1.400 ;
  END
END tt_um_tt08_aicd_playground
END LIBRARY

