* NGSPICE file created from tt_um_tt08_aicd_playground.ext - technology: sky130A

.subckt sky130_leo_ip__levelshifter_up VDDOUT VDDIN OUT IN VGND
X0 VDDIN a_373_442# a_897_442# VDDIN sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.6 as=0.3 ps=2.6 w=1 l=0.15
X1 OUT a_373_442# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.3 pd=2.6 as=0.3 ps=2.6 w=1 l=0.5
X2 VDDIN IN a_373_442# VDDIN sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.6 as=0.3 ps=2.6 w=1 l=0.15
X3 a_897_442# a_373_442# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.126 ps=1.44 w=0.42 l=0.15
X4 VDDOUT OUT a_1778_346# VDDOUT sky130_fd_pr__pfet_g5v0d10v5 ad=0.126 pd=1.44 as=0.126 ps=1.44 w=0.42 l=0.5
X5 a_1778_346# a_897_442# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.3 pd=2.6 as=0.3 ps=2.6 w=1 l=0.5
X6 VDDOUT a_1778_346# OUT VDDOUT sky130_fd_pr__pfet_g5v0d10v5 ad=0.126 pd=1.44 as=0.126 ps=1.44 w=0.42 l=0.5
X7 a_373_442# IN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.126 ps=1.44 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hvl__buf_4 VGND VNB VPWR VPB X A
X0 a_149_81# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.21 ps=1.78 w=1.5 l=0.5
X1 VGND a_149_81# X VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X2 X a_149_81# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.21375 ps=2.07 w=0.75 l=0.5
X3 X a_149_81# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X4 VPWR a_149_81# X VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X5 a_149_81# A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.105 ps=1.03 w=0.75 l=0.5
X6 VPWR a_149_81# X VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X7 X a_149_81# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.4275 ps=3.57 w=1.5 l=0.5
X8 X a_149_81# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X9 VGND a_149_81# X VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
.ends

.subckt nfet$3 a_60_n40# a_160_0# a_0_0# a_n149_n154#
X0 a_160_0# a_60_n40# a_0_0# a_n149_n154# sky130_fd_pr__nfet_g5v0d10v5 ad=0.3 pd=2.6 as=0.3 ps=2.6 w=1 l=0.5
.ends

.subckt nfet a_90_0# a_48_124# a_n123_n128# a_0_0#
X0 a_90_0# a_48_124# a_0_0# a_n123_n128# sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.126 ps=1.44 w=0.42 l=0.15
.ends

.subckt pfet$3 a_90_0# w_n184_n189# a_0_0# a_48_240#
X0 a_90_0# a_48_240# a_0_0# w_n184_n189# sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.6 as=0.3 ps=2.6 w=1 l=0.15
.ends

.subckt pfet$1 a_60_n40# w_n242_n247# a_160_0# a_0_0#
X0 a_160_0# a_60_n40# a_0_0# w_n242_n247# sky130_fd_pr__pfet_g5v0d10v5 ad=0.126 pd=1.44 as=0.126 ps=1.44 w=0.42 l=0.5
.ends

.subckt sky130_leo_ip__levelshifter_down OUT IN VGND VDDOUT
Xnfet$3_0 IN m1_306_395# VGND VGND nfet$3
Xnfet_0 OUT m1_306_395# VGND VGND nfet
Xpfet$3_0 VDDOUT VDDOUT OUT m1_306_395# pfet$3
Xpfet$1_0 IN VDDOUT VDDOUT m1_306_395# pfet$1
.ends

.subckt sky130_fd_sc_hd__and4_1 VGND VPWR VPB VNB X C A B D
X0 a_27_47# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X1 a_197_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.31245 ps=1.68 w=1 l=0.15
X3 a_303_47# C a_197_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X4 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 VPWR D a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.31245 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X6 VGND D a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.196275 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X8 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196275 ps=1.33 w=0.65 l=0.15
X9 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__mux2_1 VGND VPWR VPB VNB S A1 A0 X
X0 VPWR a_505_21# a_535_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1 a_505_21# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_218_374# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X3 VGND a_505_21# a_439_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_76_199# A0 a_218_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X5 a_505_21# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X6 a_439_47# A0 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X7 a_535_374# A1 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X8 a_76_199# A1 a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_218_47# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__dlxtp_1 VGND VPWR VPB VNB D GATE Q
X0 VPWR D a_299_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1 a_560_47# a_193_47# a_465_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.066 ps=0.745 w=0.36 l=0.15
X2 VGND a_713_21# a_659_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0936 pd=1.24 as=0.0486 ps=0.63 w=0.36 l=0.15
X3 Q a_713_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.092625 ps=0.935 w=0.65 l=0.15
X4 a_465_47# a_299_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X5 VPWR GATE a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X6 a_659_47# a_27_47# a_560_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0486 pd=0.63 as=0.0621 ps=0.705 w=0.36 l=0.15
X7 VGND a_560_47# a_713_21# VNB sky130_fd_pr__nfet_01v8 ad=0.092625 pd=0.935 as=0.169 ps=1.82 w=0.65 l=0.15
X8 VPWR a_713_21# a_644_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.07245 ps=0.765 w=0.42 l=0.15
X9 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 VPWR a_560_47# a_713_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1425 pd=1.285 as=0.26 ps=2.52 w=1 l=0.15
X11 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X12 Q a_713_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.1425 ps=1.285 w=1 l=0.15
X13 VGND D a_299_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X14 a_644_413# a_193_47# a_560_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0567 ps=0.69 w=0.42 l=0.15
X15 a_465_369# a_299_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.09575 pd=0.965 as=0.0864 ps=0.91 w=0.64 l=0.15
X16 a_560_47# a_27_47# a_465_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.09575 ps=0.965 w=0.42 l=0.15
X17 VGND GATE a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__decap_3 VPWR VGND VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=0.59
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=0.59
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VPWR VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=1.05
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=1.05
.ends

.subckt sky130_fd_sc_hd__nor3_2 VGND VPWR VPB VNB C Y A B
X0 Y C a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 a_281_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17875 ps=1.85 w=0.65 l=0.15
X6 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X10 a_281_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11 a_27_297# B a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a221o_4 VPWR VGND VPB VNB A1 B1 C1 B2 X A2
X0 VGND A2 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 VGND B2 a_1053_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2 a_804_297# B1 a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.345 pd=1.69 as=0.135 ps=1.27 w=1 l=0.15
X3 a_79_21# A1 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_445_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 a_804_297# C1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_445_297# B1 a_804_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 a_1053_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_79_21# C1 a_804_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X10 a_1053_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 a_445_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13 VGND C1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 a_804_297# B2 a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X18 a_79_21# B1 a_1053_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 a_79_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 a_445_297# B2 a_804_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.345 ps=1.69 w=1 l=0.15
X21 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 a_445_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X23 a_445_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.135 ps=1.27 w=1 l=0.15
X24 VPWR A2 a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 VPWR A1 a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1375 ps=1.275 w=1 l=0.15
X26 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X27 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfrtp_1 VGND VPWR VPB VNB Q RESET_B D CLK
X0 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X3 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X4 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X5 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X7 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X10 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X12 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X13 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X14 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X15 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X16 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X18 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X19 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X20 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X21 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X22 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X23 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X24 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X25 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X26 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X27 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_4 VGND VPWR VPB VNB X A
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X6 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X8 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X9 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_2 VPWR VGND VPB VNB X A
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a22o_1 VPWR VGND VPB VNB A1 A2 X B2 B1
X0 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X1 a_27_297# B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X2 VGND A2 a_373_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X3 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X4 a_27_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X6 a_373_47# A1 a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X7 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X8 a_109_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 a_109_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and2_1 VPWR VGND VPB VNB X B A
X0 VPWR B a_59_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 X a_59_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X2 VGND B a_145_75# VNB sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_59_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X4 X a_59_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X5 a_145_75# A a_59_75# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_2 VGND VPWR VPB VNB A X
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X1 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__and2b_1 VGND VPWR VPB VNB X A_N B
X0 VPWR B a_207_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X1 X a_207_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X2 a_297_47# a_27_413# a_207_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 X a_207_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X4 a_207_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X5 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 VGND B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X7 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__and3b_1 VGND VPWR VPB VNB A_N B X C
X0 a_109_93# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10785 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 X a_209_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X2 a_109_93# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1087 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 a_296_53# a_109_93# a_209_311# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.107825 ps=1.36 w=0.42 l=0.15
X4 VPWR C a_209_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.074375 ps=0.815 w=0.42 l=0.15
X5 a_368_53# B a_296_53# VNB sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 X a_209_311# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122275 ps=1.08 w=0.65 l=0.15
X7 a_209_311# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VPWR a_109_93# a_209_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1085 ps=1.36 w=0.42 l=0.15
X9 VGND C a_368_53# VNB sky130_fd_pr__nfet_01v8 ad=0.122275 pd=1.08 as=0.05355 ps=0.675 w=0.42 l=0.15
.ends

.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=4.73
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=4.73
.ends

.subckt sky130_fd_sc_hd__dlclkp_1 VGND VPWR VPB VNB GATE GCLK CLK
X0 a_381_369# GATE VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.09575 pd=0.965 as=0.1664 ps=1.8 w=0.64 l=0.15
X1 a_476_413# a_193_47# a_381_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.09575 ps=0.965 w=0.42 l=0.15
X2 a_957_369# a_642_307# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2032 pd=1.275 as=0.149 ps=1.325 w=0.64 l=0.15
X3 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4 a_1042_47# a_642_307# a_957_369# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 GCLK a_957_369# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.325 w=1 l=0.15
X6 VGND CLK a_1042_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0441 ps=0.63 w=0.42 l=0.15
X7 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 a_651_47# a_193_47# a_476_413# VNB sky130_fd_pr__special_nfet_01v8 ad=0.067125 pd=0.745 as=0.1192 ps=1.09 w=0.39 l=0.15
X9 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10 GCLK a_957_369# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X11 VPWR a_642_307# a_600_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X12 a_476_413# a_27_47# a_396_119# VNB sky130_fd_pr__nfet_01v8 ad=0.1192 pd=1.09 as=0.117125 ps=1.085 w=0.42 l=0.15
X13 VPWR CLK a_957_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.2032 ps=1.275 w=0.64 l=0.15
X14 a_642_307# a_476_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.118125 ps=1.04 w=0.65 l=0.15
X15 a_600_413# a_27_47# a_476_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0987 ps=0.89 w=0.42 l=0.15
X16 VPWR a_476_413# a_642_307# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.27 ps=2.54 w=1 l=0.15
X17 VGND a_642_307# a_651_47# VNB sky130_fd_pr__nfet_01v8 ad=0.118125 pd=1.04 as=0.067125 ps=0.745 w=0.42 l=0.15
X18 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X19 a_396_119# GATE VGND VNB sky130_fd_pr__nfet_01v8 ad=0.117125 pd=1.085 as=0.1281 ps=1.45 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__and3_2 VPWR VGND VPB VNB B X A C
X0 VPWR a_29_311# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_29_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.15075 ps=1.345 w=1 l=0.15
X2 VPWR A a_29_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 VGND a_29_311# X VNB sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_184_53# B a_112_53# VNB sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X5 VPWR C a_29_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15075 pd=1.345 as=0.074375 ps=0.815 w=0.42 l=0.15
X6 X a_29_311# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1304 ps=1.105 w=0.65 l=0.15
X7 a_112_53# A a_29_311# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 a_29_311# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 VGND C a_184_53# VNB sky130_fd_pr__nfet_01v8 ad=0.1304 pd=1.105 as=0.05355 ps=0.675 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o41a_4 VGND VPWR VPB VNB A1 A2 A3 A4 B1 X
X0 a_467_47# A4 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_467_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.09425 pd=0.94 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VGND A1 a_467_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.15275 ps=1.12 w=0.65 l=0.15
X3 a_467_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.09425 pd=0.94 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_467_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.15275 pd=1.12 as=0.19825 ps=1.26 w=0.65 l=0.15
X5 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.135 ps=1.27 w=1 l=0.15
X6 VPWR A1 a_1083_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 a_1083_297# A2 a_889_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VGND A3 a_467_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 a_79_21# B1 a_467_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 a_889_297# A2 a_1083_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X13 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 a_639_297# A3 a_889_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X17 VGND A2 a_467_47# VNB sky130_fd_pr__nfet_01v8 ad=0.19825 pd=1.26 as=0.09425 ps=0.94 w=0.65 l=0.15
X18 a_889_297# A3 a_639_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 a_639_297# A4 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 VPWR B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.145 ps=1.29 w=1 l=0.15
X22 VGND A4 a_467_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.09425 ps=0.94 w=0.65 l=0.15
X23 a_1083_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.49 pd=2.98 as=0.135 ps=1.27 w=1 l=0.15
X24 a_79_21# A4 a_639_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X25 a_467_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.3185 pd=2.28 as=0.08775 ps=0.92 w=0.65 l=0.15
X26 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X27 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21ai_1 VGND VPWR VPB VNB A2 A1 B1 Y
X0 Y A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X1 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X2 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X3 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X5 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__decap_6 VPWR VGND VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=1.97
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=1.97
.ends

.subckt sky130_fd_sc_hd__decap_8 VPWR VGND VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=2.89
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=2.89
.ends

.subckt sky130_fd_sc_hd__a2111o_1 VGND VPWR VPB VNB B1 X D1 A1 A2 C1
X0 VGND A2 a_660_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.082875 ps=0.905 w=0.65 l=0.15
X1 VGND C1 a_85_193# VNB sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.10075 ps=0.96 w=0.65 l=0.15
X2 a_414_297# C1 a_334_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X3 VGND a_85_193# X VNB sky130_fd_pr__nfet_01v8 ad=0.274625 pd=1.495 as=0.2145 ps=1.96 w=0.65 l=0.15
X4 a_334_297# D1 a_85_193# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X5 a_516_297# B1 a_414_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X6 a_516_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X7 a_660_47# A1 a_85_193# VNB sky130_fd_pr__nfet_01v8 ad=0.082875 pd=0.905 as=0.18525 ps=1.22 w=0.65 l=0.15
X8 a_85_193# D1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.274625 ps=1.495 w=0.65 l=0.15
X9 VPWR A1 a_516_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X10 a_85_193# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X11 VPWR a_85_193# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor2_1 VGND VPWR VPB VNB B Y A
X0 VPWR A a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_109_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor2_2 VGND VPWR VPB VNB B Y A
X0 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X5 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X7 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__dlygate4sd3_1 VGND VPWR VPB VNB A X
X0 VPWR A a_49_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 VGND a_285_47# a_391_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.5
X2 X a_391_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X3 VGND A a_49_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 VPWR a_285_47# a_391_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.5
X5 a_285_47# a_49_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X6 a_285_47# a_49_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X7 X a_391_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__diode_2 VGND VPWR VPB VNB DIODE
X0 VNB DIODE sky130_fd_pr__diode_pw2nd_05v5 perim=2.64e+06 area=4.347e+11
.ends

.subckt sky130_fd_sc_hd__and2b_2 VPWR VGND VPB VNB X B A_N
X0 VPWR a_212_413# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_297_47# a_27_413# a_212_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 X a_212_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.22895 ps=1.745 w=1 l=0.15
X3 X a_212_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.101875 ps=0.99 w=0.65 l=0.15
X4 a_212_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.07665 ps=0.785 w=0.42 l=0.15
X5 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 VPWR B a_212_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.22895 pd=1.745 as=0.0609 ps=0.71 w=0.42 l=0.15
X7 VGND B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VGND a_212_413# X VNB sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a32o_1 VGND VPWR VPB VNB X A3 B2 B1 A1 A2
X0 a_93_21# A1 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.14625 ps=1.1 w=0.65 l=0.15
X1 a_93_21# B1 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X2 a_584_47# B1 a_93_21# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X3 VPWR a_93_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2425 pd=1.485 as=0.33 ps=2.66 w=1 l=0.15
X4 VGND B2 a_584_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.06825 ps=0.86 w=0.65 l=0.15
X5 a_256_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167375 ps=1.165 w=0.65 l=0.15
X6 a_250_297# B2 a_93_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7 VGND a_93_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.167375 pd=1.165 as=0.2145 ps=1.96 w=0.65 l=0.15
X8 a_250_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.2425 ps=1.485 w=1 l=0.15
X9 VPWR A2 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X10 a_250_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X11 a_346_47# A2 a_256_47# VNB sky130_fd_pr__nfet_01v8 ad=0.14625 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o22a_1 VGND VPWR VPB VNB A2 X B1 A1 B2
X0 a_78_199# B1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1 VPWR A1 a_493_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2 a_493_297# A2 a_78_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.235 ps=1.47 w=1 l=0.15
X3 VPWR a_78_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3725 pd=1.745 as=0.28 ps=2.56 w=1 l=0.15
X4 VGND A2 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.11375 ps=1 w=0.65 l=0.15
X5 a_78_199# B2 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.235 pd=1.47 as=0.1175 ps=1.235 w=1 l=0.15
X6 a_215_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 a_215_47# B2 a_78_199# VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 a_292_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1175 pd=1.235 as=0.3725 ps=1.745 w=1 l=0.15
X9 VGND a_78_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and2_2 VPWR VGND VPB VNB A X B
X0 X a_61_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.16655 ps=1.39 w=1 l=0.15
X1 VPWR a_61_75# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.38 pd=2.76 as=0.195 ps=1.39 w=1 l=0.15
X2 VPWR B a_61_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 VGND B a_147_75# VNB sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 X a_61_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.1118 ps=1.04 w=0.65 l=0.15
X5 VGND a_61_75# X VNB sky130_fd_pr__nfet_01v8 ad=0.247 pd=2.06 as=0.12675 ps=1.04 w=0.65 l=0.15
X6 a_61_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X7 a_147_75# A a_61_75# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3_1 VPWR VGND VPB VNB A X B C
X0 X a_29_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.14825 ps=1.34 w=1 l=0.15
X1 a_111_297# C a_29_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 X a_29_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.101875 ps=0.99 w=0.65 l=0.15
X3 a_183_297# B a_111_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 VPWR A a_183_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_29_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 VGND C a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7 VGND A a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4_1 VPWR VGND VPB VNB C A X B D
X0 a_27_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_27_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_277_297# B a_205_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VPWR A a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.101875 ps=0.99 w=0.65 l=0.15
X5 a_205_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.14825 ps=1.34 w=1 l=0.15
X7 VGND C a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_109_297# D a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 VGND A a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__and3_4 VGND VPWR VPB VNB A B C X
X0 VPWR A a_94_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1975 pd=1.395 as=0.305 ps=2.61 w=1 l=0.15
X1 a_294_47# B a_185_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.128375 ps=1.045 w=0.65 l=0.15
X2 a_185_47# A a_94_47# VNB sky130_fd_pr__nfet_01v8 ad=0.128375 pd=1.045 as=0.19825 ps=1.91 w=0.65 l=0.15
X3 VPWR a_94_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X4 VGND C a_294_47# VNB sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X5 a_94_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1975 ps=1.395 w=1 l=0.15
X6 X a_94_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X7 X a_94_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X8 VPWR C a_94_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X9 X a_94_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X10 VGND a_94_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X11 VPWR a_94_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 VGND a_94_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X13 X a_94_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__or2_1 VGND VPWR VPB VNB A X B
X0 VGND A a_68_297# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_68_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 X a_68_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X3 VPWR A a_150_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 X a_68_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X5 a_150_297# B a_68_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__xnor2_1 VGND VPWR VPB VNB B Y A
X0 a_377_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.365 ps=1.73 w=1 l=0.15
X1 a_47_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3 ps=2.6 w=1 l=0.15
X2 a_129_47# B a_47_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_285_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4 Y a_47_47# a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VGND A a_129_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.06825 ps=0.86 w=0.65 l=0.15
X6 VPWR A a_47_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.365 pd=1.73 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR a_47_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.165 ps=1.33 w=1 l=0.15
X8 Y B a_377_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o2111a_1 VPWR VGND VPB VNB X D1 C1 B1 A2 A1
X0 a_676_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.2125 ps=1.425 w=1 l=0.15
X1 a_512_47# B1 a_409_47# VNB sky130_fd_pr__nfet_01v8 ad=0.19825 pd=1.26 as=0.118625 ps=1.015 w=0.65 l=0.15
X2 a_306_47# D1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.118625 pd=1.015 as=0.19825 ps=1.91 w=0.65 l=0.15
X3 VGND A2 a_512_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.19825 ps=1.26 w=0.65 l=0.15
X4 VPWR C1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.2175 ps=1.435 w=1 l=0.15
X5 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2125 pd=1.425 as=0.305 ps=1.61 w=1 l=0.15
X6 VPWR A1 a_676_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.105 ps=1.21 w=1 l=0.15
X7 a_512_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 a_409_47# C1 a_306_47# VNB sky130_fd_pr__nfet_01v8 ad=0.118625 pd=1.015 as=0.118625 ps=1.015 w=0.65 l=0.15
X9 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3825 pd=1.765 as=0.26 ps=2.52 w=1 l=0.15
X10 a_79_21# D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2175 pd=1.435 as=0.3825 ps=1.765 w=1 l=0.15
X11 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4b_4 VGND VPWR VPB VNB D_N B C A X
X0 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 VGND a_215_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VPWR a_215_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_109_93# D_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10785 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 a_215_297# a_109_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.16535 ps=1.82 w=0.65 l=0.15
X5 VGND C a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1235 ps=1.03 w=0.65 l=0.15
X6 VGND A a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X8 a_215_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_109_93# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X10 VPWR A a_487_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.135 ps=1.27 w=1 l=0.15
X11 VGND a_215_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 a_487_297# B a_403_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 a_403_297# C a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X14 VPWR a_215_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X15 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1235 ps=1.03 w=0.65 l=0.15
X16 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 a_297_297# a_109_93# a_215_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3b_4 VGND VPWR VPB VNB A B C_N X
X0 a_176_21# a_27_47# a_626_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X1 a_626_297# B a_542_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR C_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 VGND a_176_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_542_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR a_176_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 X a_176_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 X a_176_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X8 X a_176_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_176_21# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 VPWR a_176_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 X a_176_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X12 a_176_21# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X13 VGND a_176_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 VGND B a_176_21# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 VGND C_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__xor2_1 VPWR VGND VPB VNB B X A
X0 X a_35_297# a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X1 X B a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_35_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_117_297# B a_35_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 VPWR B a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND A a_35_297# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25025 ps=1.42 w=0.65 l=0.15
X7 a_285_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR A a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a22oi_1 VPWR VGND VPB VNB B1 A1 B2 A2 Y
X0 Y B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X1 Y B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.135 ps=1.27 w=1 l=0.15
X3 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 a_381_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X5 a_109_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 a_109_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X7 VGND A2 a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.234 pd=2.02 as=0.06825 ps=0.86 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o221ai_1 VGND VPWR VPB VNB A2 Y B1 C1 A1 B2
X0 a_109_47# B1 a_213_123# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1652 ps=1.82 w=0.65 l=0.15
X1 Y B2 a_295_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.12 ps=1.24 w=1 l=0.15
X2 VPWR A1 a_493_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3 a_213_123# B2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_295_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.12 pd=1.24 as=0.38 ps=1.76 w=1 l=0.15
X5 a_493_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.225 ps=1.45 w=1 l=0.15
X6 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.38 pd=1.76 as=0.28 ps=2.56 w=1 l=0.15
X7 VGND A2 a_213_123# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.117 ps=1.01 w=0.65 l=0.15
X8 a_213_123# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_109_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.1654 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfrtp_2 VGND VPWR VPB VNB Q RESET_B D CLK
X0 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X4 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X5 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X7 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X8 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X9 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X10 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X11 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X12 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X14 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X15 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X16 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X17 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X18 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X19 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X20 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X21 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X22 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X23 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X24 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X25 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X26 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X27 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X28 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X29 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21oi_1 VPWR VGND VPB VNB A1 B1 Y A2
X0 a_199_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.095875 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X1 a_113_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1475 ps=1.295 w=1 l=0.15
X2 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X3 VPWR A1 a_113_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.14 ps=1.28 w=1 l=0.15
X4 a_113_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X5 VGND A2 a_199_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.095875 ps=0.945 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o32a_1 VPWR VGND VPB VNB X A3 A1 A2 B1 B2
X0 a_77_199# B2 a_227_47# VNB sky130_fd_pr__nfet_01v8 ad=0.13325 pd=1.06 as=0.12675 ps=1.04 w=0.65 l=0.15
X1 a_323_297# A2 a_227_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.165 ps=1.33 w=1 l=0.15
X2 a_227_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3 a_227_47# B1 a_77_199# VNB sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.13325 ps=1.06 w=0.65 l=0.15
X4 VGND a_77_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5 VPWR B1 a_539_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.205 ps=1.41 w=1 l=0.15
X6 a_227_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X7 VPWR a_77_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.335 ps=2.67 w=1 l=0.15
X8 a_77_199# A3 a_323_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X9 VGND A2 a_227_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.10725 ps=0.98 w=0.65 l=0.15
X10 a_227_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 a_539_297# B2 a_77_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=1.41 as=0.195 ps=1.39 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand2_1 VGND VPWR VPB VNB Y B A
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A a_113_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_113_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o311a_1 VGND VPWR VPB VNB X A1 A2 A3 B1 C1
X0 a_585_47# B1 a_266_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.118625 ps=1.015 w=0.65 l=0.15
X1 VGND A2 a_266_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1365 pd=1.07 as=0.117 ps=1.01 w=0.65 l=0.15
X2 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3125 pd=1.625 as=0.26 ps=2.52 w=1 l=0.15
X3 a_81_21# C1 a_585_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X4 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.203125 pd=1.275 as=0.169 ps=1.82 w=0.65 l=0.15
X5 a_266_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.3125 ps=1.625 w=1 l=0.15
X6 a_368_297# A2 a_266_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.18 ps=1.36 w=1 l=0.15
X7 a_266_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.118625 pd=1.015 as=0.1365 ps=1.07 w=0.65 l=0.15
X8 a_266_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.203125 ps=1.275 w=0.65 l=0.15
X9 a_81_21# A3 a_368_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.21 ps=1.42 w=1 l=0.15
X10 a_81_21# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15 ps=1.3 w=1 l=0.15
X11 VPWR B1 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.1375 ps=1.275 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21o_2 VGND VPWR VPB VNB X B1 A1 A2
X0 VPWR a_80_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1 X a_80_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2 VGND a_80_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.1105 pd=0.99 as=0.091 ps=0.93 w=0.65 l=0.15
X3 a_386_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X4 X a_80_199# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X5 a_80_199# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1625 pd=1.15 as=0.1105 ps=0.99 w=0.65 l=0.15
X6 a_386_297# B1 a_80_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X7 a_458_47# A1 a_80_199# VNB sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.1625 ps=1.15 w=0.65 l=0.15
X8 VPWR A1 a_386_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.14 ps=1.28 w=1 l=0.15
X9 VGND A2 a_458_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.1235 ps=1.03 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o31a_1 VGND VPWR VPB VNB X A2 B1 A1 A3
X0 a_103_199# B1 a_253_47# VNB sky130_fd_pr__nfet_01v8 ad=0.2015 pd=1.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X1 VPWR a_103_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.36 ps=2.72 w=1 l=0.15
X2 a_337_297# A2 a_253_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3 a_103_199# A3 a_337_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2125 pd=1.425 as=0.165 ps=1.33 w=1 l=0.15
X4 a_253_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.195 ps=1.39 w=1 l=0.15
X5 VPWR B1 a_103_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.345 pd=2.69 as=0.2125 ps=1.425 w=1 l=0.15
X6 VGND a_103_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.234 ps=2.02 w=0.65 l=0.15
X7 a_253_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12675 ps=1.04 w=0.65 l=0.15
X8 a_253_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X9 VGND A2 a_253_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__conb_1 VGND VPWR VPB VNB LO HI
X0 VPWR HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1 LO VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
.ends

.subckt sky130_fd_sc_hd__o211a_1 VGND VPWR VPB VNB C1 B1 A2 A1 X
X0 VGND A1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1 a_510_47# B1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.143 ps=1.09 w=0.65 l=0.15
X2 a_79_21# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.175 ps=1.35 w=1 l=0.15
X3 VPWR B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.22 ps=1.44 w=1 l=0.15
X4 a_79_21# A2 a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.1625 ps=1.325 w=1 l=0.15
X5 a_297_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X6 a_79_21# C1 a_510_47# VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.11375 ps=1 w=0.65 l=0.15
X7 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X8 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X9 a_215_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.105625 ps=0.975 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a2bb2o_1 VGND VPWR VPB VNB B1 A1_N A2_N X B2
X0 a_226_47# A2_N a_226_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0441 ps=0.63 w=0.42 l=0.15
X1 a_489_413# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 a_226_297# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.16675 ps=1.435 w=0.42 l=0.15
X3 VPWR B2 a_489_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 a_489_413# a_226_47# a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 a_76_199# a_226_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1386 ps=1.08 w=0.42 l=0.15
X6 VGND B1 a_556_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 a_556_47# B2 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VGND A2_N a_226_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1386 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 a_226_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1201 ps=1.085 w=0.42 l=0.15
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16675 pd=1.435 as=0.26 ps=2.52 w=1 l=0.15
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.1201 pd=1.085 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21bo_1 VGND VPWR VPB VNB X A1 B1_N A2
X0 a_298_297# a_27_413# a_215_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1 a_215_297# a_27_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1359 ps=1.1 w=0.65 l=0.15
X2 a_298_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.258375 ps=1.445 w=0.65 l=0.15
X4 VPWR B1_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X6 a_382_47# A1 a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VGND B1_N a_27_413# VNB sky130_fd_pr__nfet_01v8 ad=0.1359 pd=1.1 as=0.1113 ps=1.37 w=0.42 l=0.15
X8 VPWR A1 a_298_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X9 VGND A2 a_382_47# VNB sky130_fd_pr__nfet_01v8 ad=0.258375 pd=1.445 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__inv_2 VPWR VGND VPB VNB A Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o2bb2a_1 VPWR VGND VPB VNB A1_N X A2_N B2 B1
X0 a_206_369# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.14575 ps=1.335 w=0.42 l=0.15
X1 a_206_369# A2_N a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06615 ps=0.735 w=0.42 l=0.15
X2 VGND B2 a_489_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_585_369# B2 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0672 ps=0.74 w=0.42 l=0.15
X4 a_489_47# a_206_369# a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 a_489_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 VPWR A2_N a_206_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.20925 pd=1.345 as=0.129 ps=1.18 w=0.42 l=0.15
X7 a_76_199# a_206_369# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.20925 ps=1.345 w=0.42 l=0.15
X8 a_205_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06615 pd=0.735 as=0.098625 ps=0.98 w=0.42 l=0.15
X9 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.26 ps=2.52 w=1 l=0.15
X10 VPWR B1 a_585_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.098625 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a211o_1 VGND VPWR VPB VNB X A2 B1 A1 C1
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X1 a_80_21# C1 a_472_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X2 VPWR A2 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.17225 ps=1.83 w=0.65 l=0.15
X5 a_300_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X6 a_217_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7 a_80_21# A1 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X8 a_472_297# B1 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X9 a_80_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor4_1 VGND VPWR VPB VNB D C Y A B
X0 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.089375 ps=0.925 w=0.65 l=0.15
X1 a_191_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.13 ps=1.26 w=1 l=0.15
X2 VPWR A a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.118625 ps=1.015 w=0.65 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 a_297_297# B a_191_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X6 a_109_297# D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.13 pd=1.26 as=0.26 ps=2.52 w=1 l=0.15
X7 Y D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.118625 pd=1.015 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4b_1 VPWR VGND VPB VNB B D_N A X C
X0 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X1 a_109_53# D_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_215_297# a_109_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.101875 ps=0.99 w=0.65 l=0.15
X4 a_392_297# C a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.04515 pd=0.635 as=0.06825 ps=0.745 w=0.42 l=0.15
X5 a_465_297# B a_392_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06405 pd=0.725 as=0.04515 ps=0.635 w=0.42 l=0.15
X6 a_215_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 VPWR A a_465_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06405 ps=0.725 w=0.42 l=0.15
X8 a_297_297# a_109_53# a_215_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 a_109_53# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X10 VGND C a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06405 ps=0.725 w=0.42 l=0.15
X11 VGND A a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_8 VGND VPWR VPB VNB X A
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.1134 pd=1.38 as=0.0588 ps=0.7 w=0.42 l=0.15
X10 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X11 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X14 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X16 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X17 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X18 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X19 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21o_1 VPWR VGND VPB VNB A2 A1 B1 X
X0 a_81_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X1 a_299_297# B1 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X2 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3 VPWR A1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X4 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X5 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X6 a_299_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7 a_384_47# A1 a_81_21# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__inv_8 VGND VPWR VPB VNB A Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3b_1 VGND VPWR VPB VNB A C_N X B
X0 a_109_93# C_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 a_215_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 VGND a_109_93# a_215_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 VGND A a_215_53# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 VPWR A a_369_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06825 ps=0.745 w=0.42 l=0.15
X5 a_369_297# B a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 X a_215_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X7 a_297_297# a_109_93# a_215_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 a_109_93# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 X a_215_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.10025 ps=0.985 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand2b_2 VGND VPWR VPB VNB B Y A_N
X0 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.335 ps=1.67 w=1 l=0.15
X1 VGND A_N a_27_93# VNB sky130_fd_pr__nfet_01v8 ad=0.194 pd=1.95 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 VGND B a_229_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 Y a_27_93# a_229_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4 a_229_47# a_27_93# Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y a_27_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.1468 ps=1.34 w=1 l=0.15
X6 VPWR a_27_93# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.335 pd=1.67 as=0.165 ps=1.33 w=1 l=0.15
X7 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.135 ps=1.27 w=1 l=0.15
X8 a_229_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VPWR A_N a_27_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1468 pd=1.34 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a221o_1 VPWR VGND VPB VNB X B1 A1 B2 A2 C1
X0 a_465_47# A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X2 a_109_297# B1 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X5 a_205_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X6 VPWR A2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X7 a_193_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X8 a_27_47# B1 a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X9 a_109_297# C1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10 VGND C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X11 VGND A2 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand3_1 VGND VPWR VPB VNB Y A C B
X0 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X2 a_193_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 Y A a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X4 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5 a_109_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor3b_4 VGND VPWR VPB VNB A C_N B Y
X0 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 VPWR A a_197_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_555_297# a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 a_197_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VGND a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 a_197_297# B a_555_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8 VGND a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VGND C_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X12 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 Y a_27_47# a_555_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 Y a_27_47# a_555_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VPWR C_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X16 a_555_297# a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 a_555_297# B a_197_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 a_197_297# B a_555_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 a_555_297# B a_197_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X22 VPWR A a_197_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X23 a_197_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25675 ps=1.44 w=0.65 l=0.15
X25 Y a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__dlxtn_1 VGND VPWR VPB VNB D GATE_N Q
X0 VPWR D a_299_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1 a_560_47# a_27_47# a_465_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.054 pd=0.66 as=0.066 ps=0.745 w=0.36 l=0.15
X2 a_465_47# a_299_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 VPWR GATE_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4 VGND a_560_47# a_715_21# VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X5 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 VPWR a_560_47# a_715_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X7 a_650_47# a_193_47# a_560_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.054 ps=0.66 w=0.36 l=0.15
X8 Q a_715_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X9 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10 VPWR a_715_21# a_644_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07455 ps=0.775 w=0.42 l=0.15
X11 VGND D a_299_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X12 Q a_715_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X13 a_644_413# a_27_47# a_560_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07455 pd=0.775 as=0.0567 ps=0.69 w=0.42 l=0.15
X14 a_465_369# a_299_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.09575 pd=0.965 as=0.0864 ps=0.91 w=0.64 l=0.15
X15 a_560_47# a_193_47# a_465_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.09575 ps=0.965 w=0.42 l=0.15
X16 VGND GATE_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X17 VGND a_715_21# a_650_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfxtp_1 VPWR VGND VPB VNB Q CLK D
X0 Q a_1059_315# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_891_413# a_193_47# a_634_159# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2 a_561_413# a_27_47# a_466_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X3 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4 Q a_1059_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 VGND a_634_159# a_592_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X7 VPWR a_891_413# a_1059_315# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X8 a_466_413# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X9 VPWR a_634_159# a_561_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X10 a_634_159# a_466_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X11 a_634_159# a_466_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X12 a_975_413# a_193_47# a_891_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 VGND a_1059_315# a_1017_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X14 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X15 a_891_413# a_27_47# a_634_159# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X16 a_592_47# a_193_47# a_466_413# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X17 VPWR a_1059_315# a_975_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X18 a_1017_47# a_27_47# a_891_413# VNB sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X19 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X20 a_466_413# a_27_47# a_381_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X21 VGND a_891_413# a_1059_315# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X22 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X23 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand2_2 VGND VPWR VPB VNB Y A B
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__inv_16 VGND VPWR VPB VNB Y A
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X17 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X22 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X26 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X28 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X29 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X30 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X31 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21a_1 VGND VPWR VPB VNB X A1 B1 A2
X0 VPWR A1 a_382_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1525 ps=1.305 w=1 l=0.15
X1 a_297_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X2 a_297_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VGND A2 a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3275 pd=1.655 as=0.28 ps=2.56 w=1 l=0.15
X5 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.3275 ps=1.655 w=1 l=0.15
X6 a_382_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.195 ps=1.39 w=1 l=0.15
X7 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor3b_2 VGND VPWR VPB VNB C_N Y A B
X0 a_281_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND a_531_21# Y VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 VPWR C_N a_531_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X7 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X9 a_281_297# a_531_21# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X10 Y a_531_21# a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X11 VGND C_N a_531_21# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X12 a_27_297# B a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X13 Y a_531_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o22ai_1 VGND VPWR VPB VNB A2 B1 Y A1 B2
X0 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X1 a_27_47# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.092625 ps=0.935 w=0.65 l=0.15
X2 VPWR A1 a_307_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.105 ps=1.21 w=1 l=0.15
X3 a_307_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.2325 ps=1.465 w=1 l=0.15
X4 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2325 pd=1.465 as=0.1125 ps=1.225 w=1 l=0.15
X6 a_109_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1125 pd=1.225 as=0.26 ps=2.52 w=1 l=0.15
X7 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.092625 pd=0.935 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_1 VGND VPWR VPB VNB X A
X0 VPWR a_75_212# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1 a_75_212# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 a_75_212# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3 VGND a_75_212# X VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand3_2 VGND VPWR VPB VNB A Y B C
X0 VGND C a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.2015 pd=1.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 a_277_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_27_47# B a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.31 pd=2.62 as=0.135 ps=1.27 w=1 l=0.15
X8 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 a_277_47# B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3_2 VGND VPWR VPB VNB A B X C
X0 VPWR a_30_53# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.315 pd=2.63 as=0.135 ps=1.27 w=1 l=0.15
X1 VGND a_30_53# X VNB sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 X a_30_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14825 ps=1.34 w=1 l=0.15
X3 a_112_297# C a_30_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 X a_30_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.101875 ps=0.99 w=0.65 l=0.15
X5 VGND A a_30_53# VNB sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 a_30_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 VGND C a_30_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 a_184_297# B a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X9 VPWR A a_184_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3b_2 VPWR VGND VPB VNB A B C_N X
X0 a_388_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.14825 ps=1.34 w=0.42 l=0.15
X1 VPWR C_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 VGND a_176_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 X a_176_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X4 VPWR a_176_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND B a_176_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 X a_176_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X7 a_176_21# a_27_47# a_472_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 a_472_297# B a_388_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 a_176_21# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.101875 ps=0.99 w=0.42 l=0.15
X10 a_176_21# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 VGND C_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4_2 VPWR VGND VPB VNB C A X B D
X0 a_27_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_27_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_277_297# B a_205_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VPWR A a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.101875 ps=0.99 w=0.65 l=0.15
X5 a_205_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 VPWR a_27_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND a_27_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.19825 pd=1.91 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14825 ps=1.34 w=1 l=0.15
X9 VGND C a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_109_297# D a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X11 VGND A a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a211oi_1 VPWR VGND VPB VNB A1 C1 B1 Y A2
X0 a_56_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VPWR A2 a_56_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
X3 a_139_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.2665 ps=2.12 w=0.65 l=0.15
X4 a_311_297# B1 a_56_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X5 Y C1 a_311_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X6 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X7 Y A1 a_139_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_16 VGND VPWR VPB VNB X A
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X6 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X7 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X14 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X16 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X17 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X18 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X19 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X20 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X21 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X22 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X23 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X24 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X25 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X26 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X27 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X28 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X29 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X30 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X31 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X32 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X33 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X34 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X35 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X36 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X37 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X38 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X39 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand2b_1 VGND VPWR VPB VNB Y A_N B
X0 VGND A_N a_27_93# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 Y a_27_93# a_206_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_206_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X3 VPWR a_27_93# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X4 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X5 VPWR A_N a_27_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_1 VGND VPWR VPB VNB X A
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkinv_16 VGND VPWR VPB VNB Y A
X0 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.14 ps=1.28 w=1 l=0.15
X3 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.2175 ps=1.435 w=1 l=0.15
X13 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.06615 pd=0.735 as=0.0588 ps=0.7 w=0.42 l=0.15
X14 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.275 ps=2.55 w=1 l=0.15
X15 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X16 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X17 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X18 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X19 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X20 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X21 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X22 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X23 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X24 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2175 pd=1.435 as=0.1575 ps=1.315 w=1 l=0.15
X25 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X26 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X27 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X28 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X29 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X30 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X31 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X32 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X33 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X34 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.09135 pd=0.855 as=0.06615 ps=0.735 w=0.42 l=0.15
X35 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X36 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X37 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X38 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X39 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.09135 ps=0.855 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o41ai_2 VGND VPWR VPB VNB A1 A2 A3 A4 Y B1
X0 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 VGND A4 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X4 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 a_299_297# A3 a_549_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X9 a_549_297# A3 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 a_299_297# A4 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 Y A4 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12 a_743_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X13 VPWR A1 a_743_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 a_743_297# A2 a_549_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 a_27_47# A4 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X16 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X17 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 a_549_297# A2 a_743_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X19 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkinv_1 VGND VPWR VPB VNB Y A
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.11 as=0.2184 ps=2.2 w=0.84 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.1197 pd=1.41 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2352 pd=2.24 as=0.1134 ps=1.11 w=0.84 l=0.15
.ends

.subckt sky130_fd_sc_hd__dlymetal6s2s_1 VPWR VGND VPB VNB A X
X0 a_558_47# a_381_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X1 VGND X a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_841_47# a_664_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X3 VPWR A a_62_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 VGND A a_62_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 a_558_47# a_381_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X6 X a_62_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X7 VPWR X a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 a_841_47# a_664_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X9 X a_62_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X10 VPWR a_558_47# a_664_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X11 VGND a_558_47# a_664_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21boi_1 VPWR VGND VPB VNB Y A1 B1_N A2
X0 a_300_297# a_27_413# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X2 VPWR B1_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.1113 ps=1.37 w=0.42 l=0.15
X3 Y a_27_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.101875 ps=0.99 w=0.65 l=0.15
X4 VPWR A1 a_300_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5 a_384_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.143 ps=1.09 w=0.65 l=0.15
X6 VGND B1_N a_27_413# VNB sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.1113 ps=1.37 w=0.42 l=0.15
X7 a_300_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__inv_12 VGND VPWR VPB VNB A Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.515 pd=3.03 as=0.135 ps=1.27 w=1 l=0.15
X4 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.33475 pd=2.33 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X14 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfrtp_4 VGND VPWR VPB VNB Q RESET_B D CLK
X0 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X3 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X4 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X5 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X12 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X14 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X15 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X16 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X17 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X18 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X19 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X20 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X21 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X22 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X23 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X24 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X25 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X26 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X27 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X28 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X29 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X30 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X31 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X32 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X33 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and3b_2 VGND VPWR VPB VNB B X A_N C
X0 a_109_53# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 X a_215_311# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12715 ps=1.095 w=0.65 l=0.15
X2 a_109_53# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 VGND C a_373_53# VNB sky130_fd_pr__nfet_01v8 ad=0.12715 pd=1.095 as=0.05355 ps=0.675 w=0.42 l=0.15
X4 VGND a_215_311# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VPWR C a_215_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.074375 ps=0.815 w=0.42 l=0.15
X6 VPWR a_215_311# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7 X a_215_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X8 a_301_53# a_109_53# a_215_311# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 a_215_311# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 a_373_53# B a_301_53# VNB sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X11 VPWR a_109_53# a_215_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a31o_1 VGND VPWR VPB VNB A2 B1 A1 A3 X
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X1 a_209_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X2 a_303_47# A2 a_209_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X3 a_209_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X5 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X6 a_80_21# A1 a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X7 VPWR A2 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X8 a_80_21# B1 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X9 a_209_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4_4 VPWR VGND VPB VNB B C A D X
X0 VPWR A a_304_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.135 ps=1.27 w=1 l=0.15
X1 a_304_297# B a_220_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND C a_32_297# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1235 ps=1.03 w=0.65 l=0.15
X3 a_220_297# C a_114_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X4 a_32_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.169 ps=1.82 w=0.65 l=0.15
X5 a_32_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VPWR a_32_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X7 X a_32_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VGND A a_32_297# VNB sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VPWR a_32_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 X a_32_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1235 ps=1.03 w=0.65 l=0.15
X11 X a_32_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 X a_32_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X13 a_114_297# D a_32_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.26 ps=2.52 w=1 l=0.15
X14 VGND a_32_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 VGND a_32_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkinvlp_4 VPWR VGND VPB VNB A Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.25
X1 VGND A a_268_47# VNB sky130_fd_pr__nfet_01v8 ad=0.14575 pd=1.63 as=0.05775 ps=0.76 w=0.55 l=0.15
X2 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.25
X3 Y A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.077 pd=0.83 as=0.05775 ps=0.76 w=0.55 l=0.15
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.25
X5 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.76 as=0.14575 ps=1.63 w=0.55 l=0.15
X6 a_268_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.76 as=0.077 ps=0.83 w=0.55 l=0.15
X7 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.25
.ends

.subckt sky130_fd_sc_hd__o221a_1 VGND VPWR VPB VNB A2 X B1 C1 A1 B2
X0 a_240_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1 X a_51_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VGND A1 a_240_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 a_51_297# B2 a_245_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.4125 pd=1.825 as=0.105 ps=1.21 w=1 l=0.15
X4 a_149_47# C1 a_51_297# VNB sky130_fd_pr__nfet_01v8 ad=0.099125 pd=0.955 as=0.2015 ps=1.92 w=0.65 l=0.15
X5 a_240_47# B1 a_149_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.099125 ps=0.955 w=0.65 l=0.15
X6 VPWR A1 a_512_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X7 X a_51_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.165 ps=1.33 w=1 l=0.15
X8 a_149_47# B2 a_240_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_245_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X10 VPWR C1 a_51_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.34 ps=2.68 w=1 l=0.15
X11 a_512_297# A2 a_51_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.4125 ps=1.825 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o211ai_1 VGND VPWR VPB VNB A1 A2 Y C1 B1
X0 a_110_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.265 ps=2.53 w=1 l=0.15
X1 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.17225 ps=1.83 w=0.65 l=0.15
X2 Y A2 a_110_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X3 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X4 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X5 a_326_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.12675 ps=1.04 w=0.65 l=0.15
X6 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.635 pd=3.27 as=0.195 ps=1.39 w=1 l=0.15
X7 Y C1 a_326_47# VNB sky130_fd_pr__nfet_01v8 ad=0.39325 pd=2.51 as=0.06825 ps=0.86 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or2_2 VPWR VGND VPB VNB B X A
X0 a_121_297# B a_39_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 X a_39_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10675 ps=1.005 w=0.65 l=0.15
X2 VPWR a_39_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 X a_39_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.15575 ps=1.355 w=1 l=0.15
X4 VGND a_39_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VPWR A a_121_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15575 pd=1.355 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 VGND A a_39_297# VNB sky130_fd_pr__nfet_01v8 ad=0.10675 pd=1.005 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 a_39_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3_4 VPWR VGND VPB VNB A X B C
X0 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.26 ps=1.45 w=0.65 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.4 ps=1.8 w=1 l=0.15
X2 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.20475 pd=1.93 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 VPWR A a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.4 pd=1.8 as=0.135 ps=1.27 w=1 l=0.15
X5 a_193_297# B a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.135 ps=1.27 w=1 l=0.15
X8 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 a_109_297# C a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13 VGND C a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21bai_1 VPWR VGND VPB VNB A1 Y B1_N A2
X0 a_388_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1275 pd=1.255 as=0.1525 ps=1.305 w=1 l=0.15
X1 a_105_352# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_297_47# a_105_352# Y VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_297_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 VPWR A1 a_388_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.1275 ps=1.255 w=1 l=0.15
X5 VGND A2 a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X6 VPWR B1_N a_105_352# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.17825 pd=1.4 as=0.1092 ps=1.36 w=0.42 l=0.15
X7 Y a_105_352# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.17825 ps=1.4 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o211ai_4 VGND VPWR VPB VNB A1 B1 A2 C1 Y
X0 VPWR A1 a_110_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 Y A2 a_110_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 a_806_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.10075 ps=0.96 w=0.65 l=0.15
X3 a_110_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 a_110_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X5 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X6 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7 a_110_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X9 VPWR A1 a_110_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.14 ps=1.28 w=1 l=0.15
X10 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_27_47# B1 a_1314_47# VNB sky130_fd_pr__nfet_01v8 ad=0.25675 pd=2.09 as=0.104 ps=0.97 w=0.65 l=0.15
X12 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X14 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X16 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X17 Y A2 a_110_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X18 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.09425 ps=0.94 w=0.65 l=0.15
X19 Y C1 a_978_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 Y C1 a_806_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X22 a_27_47# B1 a_806_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X23 a_110_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X24 a_806_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X25 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.675 pd=3.35 as=0.135 ps=1.27 w=1 l=0.15
X26 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.09425 pd=0.94 as=0.091 ps=0.93 w=0.65 l=0.15
X27 a_978_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.091 ps=0.93 w=0.65 l=0.15
X28 a_1314_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.08775 ps=0.92 w=0.65 l=0.15
X29 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X30 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.16 ps=1.32 w=1 l=0.15
X31 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o31ai_4 VGND VPWR VPB VNB A3 A2 A1 Y B1
X0 Y A3 a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_449_297# A3 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 Y A3 a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND A1 a_31_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 Y B1 a_31_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 a_449_297# A3 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.2628 ps=2.57 w=1 l=0.15
X8 Y B1 a_31_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_31_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 a_27_297# A2 a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2605 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X11 VGND A1 a_31_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12 a_31_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X14 a_31_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 a_31_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 a_449_297# A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X20 VGND A2 a_31_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X22 VGND A2 a_31_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X23 VGND A3 a_31_47# VNB sky130_fd_pr__nfet_01v8 ad=0.222625 pd=1.335 as=0.08775 ps=0.92 w=0.65 l=0.15
X24 a_31_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.222625 ps=1.335 w=0.65 l=0.15
X25 a_27_297# A2 a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X26 VGND A3 a_31_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.08775 ps=0.92 w=0.65 l=0.15
X27 a_31_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12675 ps=1.04 w=0.65 l=0.15
X28 a_449_297# A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 a_31_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X30 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X31 a_31_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o211a_2 VPWR VGND VPB VNB C1 B1 A2 A1 X
X0 a_27_47# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3675 pd=1.735 as=0.14 ps=1.28 w=1 l=0.15
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.23075 pd=2.01 as=0.091 ps=0.93 w=0.65 l=0.15
X2 VPWR C1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3 VPWR A1 a_373_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X4 a_182_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.16535 ps=1.82 w=0.65 l=0.15
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.195 ps=1.39 w=1 l=0.15
X6 a_182_47# B1 a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.16535 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.104 ps=0.97 w=0.65 l=0.15
X8 a_373_297# A2 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.3675 ps=1.735 w=1 l=0.15
X9 a_110_47# C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X10 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X11 VGND A1 a_182_47# VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21a_2 VGND VPWR VPB VNB A1 B1 A2 X
X0 VPWR A1 a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.16 ps=1.32 w=1 l=0.15
X1 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.4 ps=1.8 w=1 l=0.15
X2 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.089375 ps=0.925 w=0.65 l=0.15
X3 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.091 ps=0.93 w=0.65 l=0.15
X4 a_470_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.14 ps=1.28 w=1 l=0.15
X5 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.4 pd=1.8 as=0.1375 ps=1.275 w=1 l=0.15
X6 a_384_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X7 a_384_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.104 ps=0.97 w=0.65 l=0.15
X8 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X9 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o31a_2 VGND VPWR VPB VNB X A1 A2 B1 A3
X0 a_108_21# B1 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0.2015 pd=1.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X1 a_346_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2 X a_108_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.26325 ps=2.11 w=0.65 l=0.15
X3 a_108_21# A3 a_430_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2125 pd=1.425 as=0.165 ps=1.33 w=1 l=0.15
X4 a_430_297# A2 a_346_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR a_108_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.175 ps=1.35 w=1 l=0.15
X6 a_346_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.195 ps=1.39 w=1 l=0.15
X7 VGND A2 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 X a_108_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.405 ps=2.81 w=1 l=0.15
X9 VPWR B1 a_108_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.2125 ps=1.425 w=1 l=0.15
X10 VGND a_108_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.11375 ps=1 w=0.65 l=0.15
X11 a_346_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12675 ps=1.04 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor3_1 VGND VPWR VPB VNB C Y A B
X0 VPWR A a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_193_297# B a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_109_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and4b_4 VGND VPWR VPB VNB X D C B A_N
X0 VPWR a_174_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3275 pd=1.655 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_174_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_815_47# B a_701_47# VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.1365 ps=1.07 w=0.65 l=0.15
X3 VPWR a_174_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR C a_174_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.135 ps=1.27 w=1 l=0.15
X5 a_174_21# a_27_47# a_815_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.143 ps=1.09 w=0.65 l=0.15
X6 X a_174_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14075 ps=1.325 w=1 l=0.15
X7 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 a_701_47# C a_617_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1365 pd=1.07 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_174_21# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3275 ps=1.655 w=1 l=0.15
X10 a_174_21# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.21 ps=1.42 w=1 l=0.15
X11 VPWR a_27_47# a_174_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.22 ps=1.44 w=1 l=0.15
X12 X a_174_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X13 X a_174_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 a_617_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.212875 ps=1.305 w=0.65 l=0.15
X15 VGND a_174_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 VGND a_174_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.212875 pd=1.305 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a32oi_4 VGND VPWR VPB VNB A3 A2 A1 B1 Y B2
X0 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X2 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3375 pd=1.675 as=0.135 ps=1.27 w=1 l=0.15
X5 a_1249_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 a_1249_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2525 pd=1.505 as=0.3375 ps=1.675 w=1 l=0.15
X12 a_803_47# A2 a_1249_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.145 ps=1.29 w=1 l=0.15
X16 a_803_47# A2 a_1249_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 Y A1 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X20 Y A1 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X21 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X22 a_1249_47# A2 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.13325 ps=1.06 w=0.65 l=0.15
X23 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 a_27_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X25 a_27_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X26 a_1249_47# A2 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X27 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.2525 ps=1.505 w=1 l=0.15
X28 a_803_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.13325 pd=1.06 as=0.08775 ps=0.92 w=0.65 l=0.15
X29 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.135 ps=1.27 w=1 l=0.15
X30 a_803_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X31 VGND B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X32 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X33 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X34 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X35 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X36 VGND A3 a_1249_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X37 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X38 VGND A3 a_1249_47# VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X39 VGND B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and3b_4 VGND VPWR VPB VNB A_N X C B
X0 a_98_199# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1491 pd=1.55 as=0.108375 ps=1.01 w=0.42 l=0.15
X1 X a_56_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2 VPWR a_56_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15825 pd=1.36 as=0.14 ps=1.28 w=1 l=0.15
X3 VGND a_56_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.108375 pd=1.01 as=0.091 ps=0.93 w=0.65 l=0.15
X4 VPWR a_98_199# a_56_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1875 pd=1.375 as=0.33 ps=2.66 w=1 l=0.15
X5 VPWR a_56_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.145 ps=1.29 w=1 l=0.15
X6 VGND a_56_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X7 a_257_47# B a_152_47# VNB sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.121875 ps=1.025 w=0.65 l=0.15
X8 X a_56_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X9 X a_56_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.1775 ps=1.355 w=1 l=0.15
X10 a_152_47# a_98_199# a_56_297# VNB sky130_fd_pr__nfet_01v8 ad=0.121875 pd=1.025 as=0.19825 ps=1.91 w=0.65 l=0.15
X11 VPWR C a_56_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.15 ps=1.3 w=1 l=0.15
X12 a_98_199# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1197 pd=1.41 as=0.15825 ps=1.36 w=0.42 l=0.15
X13 a_56_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.1875 ps=1.375 w=1 l=0.15
X14 VGND C a_257_47# VNB sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.07475 ps=0.88 w=0.65 l=0.15
X15 X a_56_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o32ai_4 VGND VPWR VPB VNB A1 A2 A3 B1 Y B2
X0 a_1224_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 VPWR A1 a_1224_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1825 ps=1.365 w=1 l=0.15
X2 a_27_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1425 pd=1.285 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_806_297# A3 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.20475 ps=1.28 w=0.65 l=0.15
X8 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.20475 pd=1.28 as=0.13975 ps=1.08 w=0.65 l=0.15
X10 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_806_297# A3 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 Y A3 a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 a_27_47# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 a_27_47# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0.092625 pd=0.935 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 Y A3 a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X19 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.118625 ps=1.015 w=0.65 l=0.15
X22 a_27_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.092625 ps=0.935 w=0.65 l=0.15
X24 a_806_297# A2 a_1224_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X25 Y B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X26 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X27 VPWR B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1425 ps=1.285 w=1 l=0.15
X28 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X29 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.13975 pd=1.08 as=0.08775 ps=0.92 w=0.65 l=0.15
X30 a_1224_297# A2 a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X31 a_1224_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.135 ps=1.27 w=1 l=0.15
X32 a_806_297# A2 a_1224_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X33 VPWR A1 a_1224_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X34 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X35 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X36 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25675 ps=1.44 w=0.65 l=0.15
X37 a_1224_297# A2 a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X38 Y B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X39 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.118625 pd=1.015 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o41a_2 VGND VPWR VPB VNB A1 A2 A3 A4 B1 X
X0 VGND A2 a_393_47# VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.11375 ps=1 w=0.65 l=0.15
X1 a_496_297# A4 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.3025 ps=1.605 w=1 l=0.15
X2 a_393_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.115375 ps=1.005 w=0.65 l=0.15
X3 VPWR A1 a_697_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.41 pd=2.82 as=0.175 ps=1.35 w=1 l=0.15
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3025 pd=1.605 as=0.305 ps=1.61 w=1 l=0.15
X7 VGND A4 a_393_47# VNB sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.118625 ps=1.015 w=0.65 l=0.15
X8 a_697_297# A2 a_597_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.175 ps=1.35 w=1 l=0.15
X9 a_393_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.2665 pd=2.12 as=0.11375 ps=1 w=0.65 l=0.15
X10 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11 a_393_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.118625 pd=1.015 as=0.208 ps=1.94 w=0.65 l=0.15
X12 a_597_297# A3 a_496_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.1775 ps=1.355 w=1 l=0.15
X13 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and4b_1 VGND VPWR VPB VNB C A_N X D B
X0 a_297_47# a_27_47# a_193_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 a_369_47# B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0441 ps=0.63 w=0.42 l=0.15
X2 VPWR D a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.06615 ps=0.735 w=0.42 l=0.15
X3 X a_193_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1034 ps=1 w=0.65 l=0.15
X4 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 VGND D a_469_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1034 pd=1 as=0.0609 ps=0.71 w=0.42 l=0.15
X6 X a_193_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X7 VPWR B a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1281 pd=1.03 as=0.0987 ps=0.89 w=0.42 l=0.15
X8 a_193_413# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.1281 ps=1.03 w=0.42 l=0.15
X9 a_193_413# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 a_469_47# C a_369_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0735 ps=0.77 w=0.42 l=0.15
X11 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o41a_1 VGND VPWR VPB VNB A1 A2 A3 A4 B1 X
X0 VGND A4 a_321_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_321_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.1235 ps=1.03 w=0.65 l=0.15
X2 a_103_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=1.52 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR a_103_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.425 ps=2.85 w=1 l=0.15
X4 VGND a_103_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.247 ps=2.06 w=0.65 l=0.15
X5 VGND A2 a_321_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X6 a_321_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.12675 ps=1.04 w=0.65 l=0.15
X7 a_511_297# A3 a_393_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.22 ps=1.44 w=1 l=0.15
X8 a_619_297# A2 a_511_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X9 a_321_47# B1 a_103_21# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10 a_393_297# A4 a_103_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.26 ps=1.52 w=1 l=0.15
X11 VPWR A1 a_619_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.195 ps=1.39 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a221oi_1 VGND VPWR VPB VNB Y C1 A1 A2 B2 B1
X0 a_465_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.099125 pd=0.955 as=0.169 ps=1.82 w=0.65 l=0.15
X1 a_109_297# B1 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_204_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.069875 pd=0.865 as=0.105625 ps=0.975 w=0.65 l=0.15
X4 VGND A2 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.19825 pd=1.91 as=0.099125 ps=0.955 w=0.65 l=0.15
X5 a_193_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.26 ps=2.52 w=1 l=0.15
X6 Y B1 a_204_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.069875 ps=0.865 w=0.65 l=0.15
X7 VPWR A2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.1525 ps=1.305 w=1 l=0.15
X8 a_109_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o32a_2 VGND VPWR VPB VNB B1 B2 A3 A2 A1 X
X0 a_429_297# A2 a_345_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.215 pd=1.43 as=0.135 ps=1.27 w=1 l=0.15
X1 VGND A2 a_345_47# VNB sky130_fd_pr__nfet_01v8 ad=0.13975 pd=1.08 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.19825 pd=1.26 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_345_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.13975 ps=1.08 w=0.65 l=0.15
X5 a_345_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.305 ps=1.61 w=1 l=0.15
X6 a_629_297# B2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR B1 a_629_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.66 as=0.19 ps=1.38 w=1 l=0.15
X8 a_79_21# B2 a_345_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_345_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.2145 pd=1.96 as=0.1235 ps=1.03 w=0.65 l=0.15
X10 a_79_21# A3 a_429_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.215 ps=1.43 w=1 l=0.15
X11 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13 a_345_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.19825 ps=1.26 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__mux2_4 VPWR VGND VPB VNB X S A0 A1
X0 a_204_297# A1 a_396_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.16 ps=1.32 w=1 l=0.15
X1 VPWR a_396_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 X a_396_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR S a_314_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 a_204_297# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.1625 ps=1.325 w=1 l=0.15
X5 a_396_47# A0 a_314_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.26 ps=2.52 w=1 l=0.15
X6 a_206_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.108875 ps=0.985 w=0.65 l=0.15
X7 X a_396_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 X a_396_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VPWR a_396_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10 a_490_47# A1 a_396_47# VNB sky130_fd_pr__nfet_01v8 ad=0.274625 pd=1.495 as=0.104 ps=0.97 w=0.65 l=0.15
X11 VGND S a_490_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.274625 ps=1.495 w=0.65 l=0.15
X12 VGND a_396_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_396_47# A0 a_206_47# VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.26 ps=1.45 w=0.65 l=0.15
X14 VGND a_396_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 VPWR S a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X16 X a_396_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 VGND S a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.108875 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o31ai_1 VPWR VGND VPB VNB Y A2 A1 A3 B1
X0 Y B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.98 as=0.19825 ps=1.26 w=0.65 l=0.15
X1 Y A3 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3925 pd=1.785 as=0.135 ps=1.27 w=1 l=0.15
X2 a_193_297# A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND A2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.3925 ps=1.785 w=1 l=0.15
X5 a_109_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.19825 pd=1.26 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 a_109_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o22a_2 VGND VPWR VPB VNB A2 X B1 A1 B2
X0 a_301_47# B2 a_81_21# VNB sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 VGND A2 a_301_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1235 ps=1.03 w=0.65 l=0.15
X2 a_383_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.39 ps=1.78 w=1 l=0.15
X3 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.39 pd=1.78 as=0.135 ps=1.27 w=1 l=0.15
X4 a_301_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 X a_81_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7 X a_81_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X8 VPWR A1 a_579_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.105 ps=1.21 w=1 l=0.15
X9 a_81_21# B1 a_301_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10 a_579_297# A2 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.235 ps=1.47 w=1 l=0.15
X11 a_81_21# B2 a_383_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.235 pd=1.47 as=0.105 ps=1.21 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__and4_2 VGND VPWR VPB VNB X C A B D
X0 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.10725 ps=0.98 w=0.65 l=0.15
X1 VGND D a_304_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17515 pd=1.265 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.27995 ps=1.615 w=1 l=0.15
X3 a_198_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.06195 ps=0.715 w=0.42 l=0.15
X4 a_27_47# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X5 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.165 ps=1.33 w=1 l=0.15
X6 a_304_47# C a_198_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X7 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07455 pd=0.775 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 VPWR D a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27995 pd=1.615 as=0.0588 ps=0.7 w=0.42 l=0.15
X9 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.17515 ps=1.265 w=0.65 l=0.15
X10 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.07455 ps=0.775 w=0.42 l=0.15
X11 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__dlxtn_2 VPWR VGND VPB VNB D GATE_N Q
X0 VPWR a_728_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 VGND a_728_21# a_663_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2 VPWR a_728_21# a_686_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VPWR GATE_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4 a_686_413# a_27_47# a_565_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.09555 ps=0.875 w=0.42 l=0.15
X5 VGND a_728_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 Q a_728_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1425 ps=1.285 w=1 l=0.15
X7 VGND a_565_413# a_728_21# VNB sky130_fd_pr__nfet_01v8 ad=0.092625 pd=0.935 as=0.169 ps=1.82 w=0.65 l=0.15
X8 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 a_663_47# a_193_47# a_565_413# VNB sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0504 ps=0.64 w=0.36 l=0.15
X10 a_469_369# a_303_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0968 pd=0.97 as=0.0864 ps=0.91 w=0.64 l=0.15
X11 VGND D a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X12 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X13 VPWR D a_303_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X14 a_565_413# a_193_47# a_469_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.09555 pd=0.875 as=0.0968 ps=0.97 w=0.42 l=0.15
X15 VPWR a_565_413# a_728_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1425 pd=1.285 as=0.26 ps=2.52 w=1 l=0.15
X16 a_469_47# a_303_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0777 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 VGND GATE_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X18 a_565_413# a_27_47# a_469_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0504 pd=0.64 as=0.0777 ps=0.81 w=0.36 l=0.15
X19 Q a_728_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.092625 ps=0.935 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor2_4 VGND VPWR VPB VNB Y A B
X0 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X6 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X11 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4bb_1 VPWR VGND VPB VNB A X B D_N C_N
X0 VGND A a_311_413# VNB sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 VPWR A a_561_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.05985 ps=0.705 w=0.42 l=0.15
X2 a_393_413# a_205_93# a_311_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1215 pd=1.33 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 VGND C_N a_27_410# VNB sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 VPWR C_N a_27_410# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1226 pd=1.32 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 X a_311_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X6 VGND a_27_410# a_311_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.05985 ps=0.705 w=0.42 l=0.15
X7 a_561_297# B a_489_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.05985 pd=0.705 as=0.0441 ps=0.63 w=0.42 l=0.15
X8 a_205_93# D_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06195 ps=0.715 w=0.42 l=0.15
X9 a_205_93# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.1226 ps=1.32 w=0.42 l=0.15
X10 a_489_297# a_27_410# a_393_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1215 ps=1.33 w=0.42 l=0.15
X11 a_311_413# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X12 a_311_413# a_205_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.05985 pd=0.705 as=0.1092 ps=1.36 w=0.42 l=0.15
X13 X a_311_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.101875 ps=0.99 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21oi_2 VGND VPWR VPB VNB B1 A2 A1 Y
X0 VGND A2 a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.06825 ps=0.86 w=0.65 l=0.15
X1 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.26 pd=2.1 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 Y A1 a_114_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X3 a_114_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.18525 ps=1.87 w=0.65 l=0.15
X4 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.135 ps=1.27 w=1 l=0.15
X5 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.15
X8 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X10 a_285_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.091 ps=0.93 w=0.65 l=0.15
X11 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o2111a_2 VGND VPWR VPB VNB D1 C1 A2 A1 B1 X
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.365 pd=1.73 as=0.14 ps=1.28 w=1 l=0.15
X1 X a_80_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2 a_80_21# D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.365 ps=1.73 w=1 l=0.15
X3 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X4 VPWR C1 a_80_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.14 ps=1.28 w=1 l=0.15
X5 X a_80_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X6 a_80_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X7 a_674_297# A2 a_80_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X8 a_386_47# D1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X9 VPWR A1 a_674_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.195 ps=1.39 w=1 l=0.15
X10 a_566_47# B1 a_458_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X11 VGND A2 a_566_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X12 a_566_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.12675 ps=1.04 w=0.65 l=0.15
X13 a_458_47# C1 a_386_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.06825 ps=0.86 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4b_2 VPWR VGND VPB VNB C A X B D_N
X0 a_176_21# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 VGND D_N a_27_53# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 VGND a_176_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 X a_176_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X4 VPWR a_176_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16835 pd=1.495 as=0.135 ps=1.27 w=1 l=0.15
X5 a_555_297# C a_483_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 a_176_21# a_27_53# a_555_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 X a_176_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1693 ps=1.5 w=1 l=0.15
X8 a_387_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.16835 ps=1.495 w=0.42 l=0.15
X9 a_483_297# B a_387_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 VGND B a_176_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X11 VGND a_27_53# a_176_21# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12 VPWR D_N a_27_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1693 pd=1.5 as=0.1092 ps=1.36 w=0.42 l=0.15
X13 a_176_21# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.10025 ps=0.985 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o32ai_2 VGND VPWR VPB VNB A1 B1 A2 A3 Y B2
X0 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25675 ps=1.44 w=0.65 l=0.15
X1 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25675 ps=1.44 w=0.65 l=0.15
X2 a_475_297# A2 a_729_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X3 a_729_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 VPWR A1 a_729_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X5 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_27_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7 a_729_297# A2 a_475_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_27_47# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_475_297# A3 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 Y A3 a_475_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X15 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.2275 pd=2 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X19 Y B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_4 VPWR VGND VPB VNB X A
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21ba_1 VGND VPWR VPB VNB B1_N A1 X A2
X0 a_222_93# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X1 VPWR A1 a_544_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.105 ps=1.21 w=1 l=0.15
X2 VGND a_79_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_222_93# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.18575 ps=1.415 w=0.42 l=0.15
X4 VGND A2 a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X5 a_448_47# a_222_93# a_79_199# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X6 a_79_199# a_222_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.3 ps=2.6 w=1 l=0.15
X7 a_544_297# A2 a_79_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X8 a_448_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VPWR a_79_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18575 pd=1.415 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__mux4_1 VGND VPWR VPB VNB S0 A1 X S1 A2 A0 A3
X0 a_277_47# a_247_21# a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 VGND S0 a_247_21# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_834_97# a_247_21# a_750_97# VNB sky130_fd_pr__nfet_01v8 ad=0.10795 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 VGND A3 a_668_97# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1079 ps=1.36 w=0.42 l=0.15
X4 a_1290_413# S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 a_834_97# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 a_750_97# S0 a_757_363# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1079 ps=1.36 w=0.42 l=0.15
X7 a_27_47# S0 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.085225 ps=0.925 w=0.42 l=0.15
X8 X a_1478_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X9 VPWR A1 a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10 VPWR S0 a_247_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1079 pd=1.36 as=0.1083 ps=1.36 w=0.42 l=0.15
X11 X a_1478_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X12 a_193_47# A0 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 a_750_97# a_1290_413# a_1478_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2688 pd=2.12 as=0.092075 ps=0.99 w=0.42 l=0.15
X14 a_1478_413# S1 a_277_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.092075 pd=0.99 as=0.1092 ps=1.36 w=0.42 l=0.15
X15 a_1290_413# S1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X16 a_277_47# a_247_21# a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0.085225 pd=0.925 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 a_750_97# S0 a_668_97# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X18 a_923_363# a_247_21# a_750_97# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.090125 pd=0.995 as=0.0567 ps=0.69 w=0.42 l=0.15
X19 a_757_363# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X20 VPWR A3 a_923_363# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.090125 ps=0.995 w=0.42 l=0.15
X21 a_277_47# a_1290_413# a_1478_413# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.151025 ps=1.285 w=0.42 l=0.15
X22 a_193_413# A0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X23 a_193_413# S0 a_277_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1079 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X24 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X25 a_1478_413# S1 a_750_97# VNB sky130_fd_pr__nfet_01v8 ad=0.151025 pd=1.285 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o22ai_4 VGND VPWR VPB VNB A1 Y A2 B1 B2
X0 a_33_47# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 VGND A1 a_33_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VGND A2 a_33_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 a_33_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_797_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 Y A2 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_797_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 Y B2 a_797_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 a_115_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VPWR B1 a_797_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 a_33_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VGND A1 a_33_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12 a_33_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_33_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 Y A2 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 a_33_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 a_797_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.16 ps=1.32 w=1 l=0.15
X17 a_115_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 VPWR A1 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 VPWR B1 a_797_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X20 VGND A2 a_33_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 a_33_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 a_797_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 VPWR A1 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.135 ps=1.27 w=1 l=0.15
X24 Y B2 a_33_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X25 Y B2 a_797_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X26 Y B1 a_33_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.104 ps=0.97 w=0.65 l=0.15
X27 Y B2 a_33_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X28 a_115_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 Y B1 a_33_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X30 a_33_47# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X31 a_115_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.29 ps=2.58 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a41o_4 VGND VPWR VPB VNB X A4 A3 A2 A1 B1
X0 a_639_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_639_47# A2 a_889_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR A3 a_467_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.385 pd=1.77 as=0.145 ps=1.29 w=1 l=0.15
X4 a_889_47# A2 a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 a_889_47# A3 a_1079_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_467_297# A4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.09425 pd=0.94 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 a_467_297# B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.135 ps=1.27 w=1 l=0.15
X13 a_467_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.135 ps=1.27 w=1 l=0.15
X14 VPWR A4 a_467_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 a_1079_47# A3 a_889_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 a_79_21# B1 a_467_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X17 a_79_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.09425 ps=0.94 w=0.65 l=0.15
X18 a_1079_47# A4 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 VPWR A2 a_467_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 a_467_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X22 a_79_21# A1 a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X23 VPWR A1 a_467_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.145 ps=1.29 w=1 l=0.15
X24 a_467_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.385 ps=1.77 w=1 l=0.15
X25 VGND A4 a_1079_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X26 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X27 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o32a_4 VGND VPWR VPB VNB X B2 A1 A2 A3 B1
X0 a_27_47# B2 a_549_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 VGND a_549_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VPWR a_549_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 a_27_297# A2 a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4 a_277_297# A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 a_549_297# B2 a_739_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.135 ps=1.27 w=1 l=0.15
X6 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 a_739_297# B2 a_549_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15 ps=1.3 w=1 l=0.15
X9 a_739_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.09425 pd=0.94 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 a_549_297# B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0975 ps=0.95 w=0.65 l=0.15
X13 a_277_297# A3 a_549_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X14 VPWR B1 a_739_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15 X a_549_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 a_27_47# B1 a_549_297# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X17 a_549_297# A3 a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X18 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.09425 ps=0.94 w=0.65 l=0.15
X19 VPWR a_549_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VGND a_549_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 X a_549_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X23 a_549_297# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X24 X a_549_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X25 X a_549_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X26 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X27 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a41oi_4 VGND VPWR VPB VNB B1 A2 A1 A4 A3 Y
X0 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.29 ps=1.58 w=1 l=0.15
X1 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.3375 ps=1.675 w=1 l=0.15
X2 Y A1 a_493_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR A4 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 Y A1 a_493_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.305 ps=1.61 w=1 l=0.15
X6 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1825 ps=1.365 w=1 l=0.15
X7 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 a_911_47# A2 a_493_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_911_47# A3 a_1269_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 VGND A4 a_1269_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 VGND A4 a_1269_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=1.58 as=0.135 ps=1.27 w=1 l=0.15
X14 a_493_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 a_493_47# A2 a_911_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 a_493_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 a_493_47# A2 a_911_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 a_911_47# A2 a_493_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X23 a_1269_47# A4 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.08775 ps=0.92 w=0.65 l=0.15
X24 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.135 ps=1.27 w=1 l=0.15
X26 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.145 ps=1.29 w=1 l=0.15
X27 a_911_47# A3 a_1269_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X28 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X29 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X30 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3375 pd=1.675 as=0.135 ps=1.27 w=1 l=0.15
X31 a_27_297# A4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X32 VPWR A4 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X33 a_1269_47# A3 a_911_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X34 a_27_297# A4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X35 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X36 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X37 a_1269_47# A3 a_911_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X38 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X39 a_1269_47# A4 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt dig_ctrl_top clk ena rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5]
+ uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7]
+ uio_oe[0] uio_oe[1] uio_oe[3] uio_oe[4] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1]
+ uio_out[2] uio_out[3] uio_out[4] uio_out[6] uio_out[7] uo_out[0] uo_out[1] uo_out[2]
+ uo_out[3] uo_out[4] uo_out[5] uo_out[6] uo_out[7] clk_o port_ms_i port_ms_o[0] port_ms_o[1]
+ port_ms_o[2] port_ms_o[3] port_ms_o[4] port_ms_o[5] port_ms_o[6] port_ms_o[7] uio_out[5]
+ ui_in[6] uio_oe[5] uio_oe[2] ui_in[7] VGND VDPWR
X_2037_ VGND VDPWR VDPWR VGND _0696_ net115 dig_ctrl_inst.latch_mem_inst.RAM\[14\]\[6\]
+ net129 net78 sky130_fd_sc_hd__and4_1
X_2106_ VGND VDPWR VDPWR VGND _0762_ _0340_ dig_ctrl_inst.cpu_inst.data\[0\] _0035_
+ sky130_fd_sc_hd__mux2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[41\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND net215 dig_ctrl_inst.latch_mem_inst.gclk\[41\] dig_ctrl_inst.latch_mem_inst.RAM\[41\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_15_Left_93 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[30\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND net234 dig_ctrl_inst.latch_mem_inst.gclk\[30\] dig_ctrl_inst.latch_mem_inst.RAM\[30\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_2_119 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_64_25 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1270_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[0\]\[3\] _1112_ net254
+ net250 sky130_fd_sc_hd__nor3_2
X_1606_ VDPWR VGND VDPWR VGND net136 net102 _1172_ _1106_ _0271_ net122 sky130_fd_sc_hd__a221o_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[56\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND net191 dig_ctrl_inst.latch_mem_inst.gclk\[56\] dig_ctrl_inst.latch_mem_inst.RAM\[56\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_38_81 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2586_ VGND VDPWR VDPWR VGND net20 net173 _0100_ clknet_leaf_6_clk sky130_fd_sc_hd__dfrtp_1
Xfanout138 VGND VDPWR VDPWR VGND net138 _1140_ sky130_fd_sc_hd__clkbuf_4
Xfanout127 VDPWR VGND VDPWR VGND net127 net131 sky130_fd_sc_hd__buf_2
X_1468_ VDPWR VGND VDPWR VGND net264 dig_ctrl_inst.spi_data_o\[3\] dig_ctrl_inst.data_out\[3\]
+ _0164_ _1113_ sky130_fd_sc_hd__a22o_1
X_1399_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[30\] _0132_ net147
+ sky130_fd_sc_hd__and2_1
Xfanout149 VDPWR VGND VDPWR VGND net149 _1081_ sky130_fd_sc_hd__buf_2
Xfanout105 VGND VDPWR VDPWR VGND _1179_ net105 sky130_fd_sc_hd__clkbuf_2
X_1537_ VGND VDPWR VDPWR VGND _0191_ net160 dig_ctrl_inst.cpu_inst.data\[2\] _0207_
+ sky130_fd_sc_hd__mux2_1
Xfanout116 VDPWR VGND VDPWR VGND net116 net118 sky130_fd_sc_hd__buf_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[45\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND net210 dig_ctrl_inst.latch_mem_inst.gclk\[45\] dig_ctrl_inst.latch_mem_inst.RAM\[45\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_64_158 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[34\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND net222 dig_ctrl_inst.latch_mem_inst.gclk\[34\] dig_ctrl_inst.latch_mem_inst.RAM\[34\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_0_Left_78 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[23\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND net238 dig_ctrl_inst.latch_mem_inst.gclk\[23\] dig_ctrl_inst.latch_mem_inst.RAM\[23\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
X_2440_ VGND VDPWR VDPWR VGND _1025_ _1022_ _1023_ sky130_fd_sc_hd__and2b_1
X_1322_ VGND VDPWR VDPWR VGND net263 net259 _1164_ dig_ctrl_inst.cpu_inst.regs\[2\]\[4\]
+ sky130_fd_sc_hd__and3b_1
X_2371_ VGND VDPWR VDPWR VGND _0991_ _1001_ net344 _0061_ sky130_fd_sc_hd__mux2_1
X_1253_ VGND VDPWR VDPWR VGND net249 dig_ctrl_inst.cpu_inst.regs\[1\]\[1\] _1095_
+ net253 sky130_fd_sc_hd__and3b_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[11\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND net183 dig_ctrl_inst.latch_mem_inst.gclk\[11\] dig_ctrl_inst.latch_mem_inst.RAM\[11\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_6_266 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_309 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2569_ VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_receiver_inst.synchronizer_spi_sclk.pipe\[0\]
+ net168 net13 clknet_leaf_4_clk sky130_fd_sc_hd__dfrtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[49\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND net198 dig_ctrl_inst.latch_mem_inst.gclk\[49\] dig_ctrl_inst.latch_mem_inst.RAM\[49\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[5\].gen_latches\[0\].p_latch VGND VDPWR VDPWR
+ VGND net237 dig_ctrl_inst.latch_mem_inst.gclk\[5\] dig_ctrl_inst.latch_mem_inst.RAM\[5\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_27_Left_105 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.genblk1\[16\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[16\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[16\]._gclk clknet_leaf_16_clk sky130_fd_sc_hd__dlclkp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[38\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND net218 dig_ctrl_inst.latch_mem_inst.gclk\[38\] dig_ctrl_inst.latch_mem_inst.RAM\[38\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_36_Left_114 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_45_Left_123 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[27\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND net231 dig_ctrl_inst.latch_mem_inst.gclk\[27\] dig_ctrl_inst.latch_mem_inst.RAM\[27\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
X_1871_ VDPWR VGND VDPWR VGND net94 _0532_ dig_ctrl_inst.latch_mem_inst.RAM\[38\]\[4\]
+ net53 sky130_fd_sc_hd__and3_2
XPHY_EDGE_ROW_54_Left_132 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1940_ VGND VDPWR VDPWR VGND _0600_ net75 dig_ctrl_inst.latch_mem_inst.RAM\[46\]\[5\]
+ net114 net52 sky130_fd_sc_hd__and4_1
XFILLER_0_16_309 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_2423_ VGND VDPWR VDPWR VGND net139 dig_ctrl_inst.cpu_inst.port_o\[5\] net327 _0101_
+ sky130_fd_sc_hd__mux2_1
X_2285_ VDPWR VGND VDPWR VGND dig_ctrl_inst.spi_data_o\[4\] _0183_ _0927_ dig_ctrl_inst.synchronizer_port_i_inst\[4\].out
+ _0824_ sky130_fd_sc_hd__a22o_1
X_1305_ VGND VDPWR VDPWR VGND _1063_ _1143_ _1144_ _1145_ _1146_ _1147_ sky130_fd_sc_hd__o41a_4
X_2354_ VGND VDPWR VDPWR VGND _0766_ net166 _0822_ _0992_ sky130_fd_sc_hd__o21ai_1
X_1236_ VGND VDPWR VDPWR VGND _1078_ net255 dig_ctrl_inst.cpu_inst.regs\[2\]\[0\]
+ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_63_Left_141 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_19_50 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_72_Left_150 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[9\].gen_latches\[1\].p_latch VGND VDPWR VDPWR
+ VGND net228 dig_ctrl_inst.latch_mem_inst.gclk\[9\] dig_ctrl_inst.latch_mem_inst.RAM\[9\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_25_128 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_25_139 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_2070_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[45\]\[7\] _0147_ _0728_
+ dig_ctrl_inst.latch_mem_inst.RAM\[5\]\[7\] _0272_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_3_Left_81 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_72_25 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1854_ VGND VDPWR VDPWR VGND _0469_ _0516_ _0492_ dig_ctrl_inst.latch_mem_inst.RAM\[9\]\[3\]
+ _1188_ _0470_ sky130_fd_sc_hd__a2111o_1
X_1785_ VDPWR VGND VDPWR VGND net95 _0448_ dig_ctrl_inst.latch_mem_inst.RAM\[38\]\[2\]
+ net57 sky130_fd_sc_hd__and3_2
X_1923_ VDPWR VGND VDPWR VGND net86 _0583_ dig_ctrl_inst.latch_mem_inst.RAM\[56\]\[5\]
+ net45 sky130_fd_sc_hd__and3_2
X_2406_ VGND VDPWR VDPWR VGND _0176_ dig_ctrl_inst.spi_data_o\[6\] dig_ctrl_inst.spi_data_o\[5\]
+ _0086_ sky130_fd_sc_hd__mux2_1
X_2268_ VGND VDPWR VDPWR VGND net150 _0798_ _0780_ _0910_ sky130_fd_sc_hd__mux2_1
X_1219_ VGND VDPWR VDPWR VGND net257 _1061_ net261 sky130_fd_sc_hd__nor2_1
X_2199_ VGND VDPWR VDPWR VGND net176 _0844_ _1060_ sky130_fd_sc_hd__nor2_2
X_2337_ VDPWR VGND VDPWR VGND dig_ctrl_inst.cpu_inst.data\[7\] _0813_ _0976_ _0227_
+ _0844_ sky130_fd_sc_hd__a22o_1
Xhold63 VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[3\]\[6\] net345 sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[3\]\[7\] net334 sky130_fd_sc_hd__dlygate4sd3_1
Xhold30 VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[3\]\[5\] net312 sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 VGND VDPWR VDPWR VGND net20 net356 sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[1\]\[2\] net323 sky130_fd_sc_hd__dlygate4sd3_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[60\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND net229 dig_ctrl_inst.latch_mem_inst.gclk\[60\] dig_ctrl_inst.latch_mem_inst.RAM\[60\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_38_253 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_5 VGND VDPWR VDPWR VGND _0379_ sky130_fd_sc_hd__diode_2
XFILLER_0_21_164 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1570_ VGND VDPWR VDPWR VGND _0235_ _0236_ _0233_ sky130_fd_sc_hd__nor2_1
X_2122_ VDPWR VGND VDPWR VGND _0768_ _0767_ _0766_ sky130_fd_sc_hd__and2b_2
X_2053_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[33\]\[7\] _0136_ _0711_
+ dig_ctrl_inst.latch_mem_inst.RAM\[36\]\[7\] _0139_ sky130_fd_sc_hd__a22o_1
X_1768_ VGND VDPWR VDPWR VGND _0431_ net78 dig_ctrl_inst.latch_mem_inst.RAM\[45\]\[2\]
+ net121 net56 sky130_fd_sc_hd__and4_1
X_1837_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[35\]\[3\] _0138_ _0499_
+ dig_ctrl_inst.latch_mem_inst.RAM\[46\]\[3\] _0148_ sky130_fd_sc_hd__a22o_1
X_1906_ VGND VDPWR VDPWR VGND _0567_ net39 dig_ctrl_inst.latch_mem_inst.RAM\[19\]\[4\]
+ _0124_ dig_ctrl_inst.latch_mem_inst.RAM\[54\]\[4\] net93 sky130_fd_sc_hd__a32o_1
X_1699_ VGND VDPWR VDPWR VGND _0360_ _0363_ _0362_ dig_ctrl_inst.latch_mem_inst.RAM\[62\]\[1\]
+ _0162_ _0361_ sky130_fd_sc_hd__a2111o_1
Xoutput20 VDPWR VGND VDPWR VGND port_ms_o[4] net20 sky130_fd_sc_hd__buf_2
Xoutput31 VDPWR VGND VDPWR VGND uo_out[6] net31 sky130_fd_sc_hd__buf_2
XFILLER_0_73_329 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
Xdig_ctrl_inst.latch_mem_inst.gen_words\[53\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND net241 dig_ctrl_inst.latch_mem_inst.gclk\[53\] dig_ctrl_inst.latch_mem_inst.RAM\[53\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
X_1622_ VDPWR VGND VDPWR VGND net81 _0287_ dig_ctrl_inst.latch_mem_inst.RAM\[26\]\[0\]
+ net66 sky130_fd_sc_hd__and3_2
XFILLER_0_1_312 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1484_ VGND VDPWR VDPWR VGND net167 dig_ctrl_inst.cpu_inst.stb_o _0173_ _1073_ _0175_
+ sky130_fd_sc_hd__o22a_1
X_1553_ VDPWR VGND VDPWR VGND net258 _0219_ net262 dig_ctrl_inst.cpu_inst.regs\[3\]\[7\]
+ sky130_fd_sc_hd__and3_2
XFILLER_0_49_337 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2036_ VDPWR VGND VDPWR VGND net129 _0695_ dig_ctrl_inst.latch_mem_inst.RAM\[4\]\[6\]
+ net98 sky130_fd_sc_hd__and3_2
X_2105_ VDPWR VGND VDPWR VGND _1055_ _0762_ _0194_ sky130_fd_sc_hd__and2_2
XFILLER_0_64_318 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[41\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND net182 dig_ctrl_inst.latch_mem_inst.gclk\[41\] dig_ctrl_inst.latch_mem_inst.RAM\[41\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[30\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND net200 dig_ctrl_inst.latch_mem_inst.gclk\[30\] dig_ctrl_inst.latch_mem_inst.RAM\[30\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[0\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[0\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[0\]._gclk clknet_leaf_14_clk sky130_fd_sc_hd__dlclkp_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[23\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[23\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[23\]._gclk clknet_leaf_13_clk sky130_fd_sc_hd__dlclkp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[57\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND net228 dig_ctrl_inst.latch_mem_inst.gclk\[57\] dig_ctrl_inst.latch_mem_inst.RAM\[57\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_73_148 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_13_52 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2585_ VGND VDPWR VDPWR VGND net19 net173 _0099_ clknet_leaf_6_clk sky130_fd_sc_hd__dfrtp_1
X_1605_ VDPWR VGND VDPWR VGND _1053_ _0270_ _0194_ sky130_fd_sc_hd__and2_2
X_1536_ VDPWR VGND VDPWR VGND dig_ctrl_inst.cpu_inst.ip\[2\] _0206_ _0185_ _0200_
+ sky130_fd_sc_hd__or3_1
Xfanout128 VGND VDPWR VDPWR VGND net131 net128 sky130_fd_sc_hd__clkbuf_2
X_1467_ VDPWR VGND VDPWR VGND net264 dig_ctrl_inst.spi_data_o\[2\] dig_ctrl_inst.data_out\[2\]
+ _0164_ _1129_ sky130_fd_sc_hd__a22o_1
Xfanout106 VDPWR VGND VDPWR VGND net106 net110 sky130_fd_sc_hd__buf_2
X_1398_ VDPWR VGND VDPWR VGND net78 _0132_ net115 net68 sky130_fd_sc_hd__and3_2
Xfanout117 VGND VDPWR VDPWR VGND net118 net117 sky130_fd_sc_hd__clkbuf_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[1\].gen_latches\[3\].p_latch VGND VDPWR VDPWR
+ VGND net215 dig_ctrl_inst.latch_mem_inst.gclk\[1\] dig_ctrl_inst.latch_mem_inst.RAM\[1\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
X_2019_ VGND VDPWR VDPWR VGND _0678_ net101 dig_ctrl_inst.latch_mem_inst.RAM\[55\]\[6\]
+ net109 net47 sky130_fd_sc_hd__and4_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[34\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND net188 dig_ctrl_inst.latch_mem_inst.gclk\[34\] dig_ctrl_inst.latch_mem_inst.RAM\[34\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[23\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND net206 dig_ctrl_inst.latch_mem_inst.gclk\[23\] dig_ctrl_inst.latch_mem_inst.RAM\[23\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[32\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[32\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[32\]._gclk sky130_fd_sc_hd__clkbuf_4
X_1321_ VDPWR VGND VDPWR VGND _1070_ _1163_ _1055_ _1162_ sky130_fd_sc_hd__and3_2
X_1252_ VGND VDPWR VDPWR VGND net253 net249 _1094_ dig_ctrl_inst.cpu_inst.regs\[2\]\[1\]
+ sky130_fd_sc_hd__and3b_1
X_2370_ VDPWR VGND VDPWR VGND _0986_ _0974_ _1001_ _0982_ _1000_ sky130_fd_sc_hd__or4_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[12\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND net219 dig_ctrl_inst.latch_mem_inst.gclk\[12\] dig_ctrl_inst.latch_mem_inst.RAM\[12\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_6_278 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_2568_ VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_receiver_inst.spi_cs_sync net170 net295
+ clknet_leaf_4_clk sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_12_Right_12 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2499_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.ip\[5\] net152 _0025_ clknet_leaf_14_clk
+ sky130_fd_sc_hd__dfrtp_1
X_1519_ VGND VDPWR VDPWR VGND _1076_ _0191_ _1062_ sky130_fd_sc_hd__nor2_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[5\].gen_latches\[4\].p_latch VGND VDPWR VDPWR
+ VGND net203 dig_ctrl_inst.latch_mem_inst.gclk\[5\] dig_ctrl_inst.latch_mem_inst.RAM\[5\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_21_Right_21 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_4_72 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_45_181 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
Xdig_ctrl_inst.latch_mem_inst.gen_words\[38\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND net181 dig_ctrl_inst.latch_mem_inst.gclk\[38\] dig_ctrl_inst.latch_mem_inst.RAM\[38\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_30_Right_30 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_29_29 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
Xdig_ctrl_inst.latch_mem_inst.gen_words\[27\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND net199 dig_ctrl_inst.latch_mem_inst.gclk\[27\] dig_ctrl_inst.latch_mem_inst.RAM\[27\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_28_104 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_1870_ VGND VDPWR VDPWR VGND _0531_ net77 dig_ctrl_inst.latch_mem_inst.RAM\[61\]\[4\]
+ net119 _0150_ sky130_fd_sc_hd__and4_1
XFILLER_0_3_204 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[16\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND net211 dig_ctrl_inst.latch_mem_inst.gclk\[16\] dig_ctrl_inst.latch_mem_inst.RAM\[16\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
X_2422_ VGND VDPWR VDPWR VGND net139 dig_ctrl_inst.cpu_inst.port_o\[4\] net356 _0100_
+ sky130_fd_sc_hd__mux2_1
X_2353_ VGND VDPWR VDPWR VGND _1068_ _0189_ _0769_ _0991_ sky130_fd_sc_hd__and3_4
X_2284_ VGND VDPWR VDPWR VGND _0924_ _0926_ _0925_ sky130_fd_sc_hd__or2_1
X_1304_ VDPWR VGND VDPWR VGND net256 _1146_ net251 dig_ctrl_inst.cpu_inst.regs\[0\]\[5\]
+ sky130_fd_sc_hd__or3_1
X_1235_ VDPWR VGND VDPWR VGND net255 _1077_ dig_ctrl_inst.cpu_inst.regs\[3\]\[0\]
+ net251 sky130_fd_sc_hd__and3_2
X_1999_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[13\]\[6\] _0117_ _0658_
+ dig_ctrl_inst.latch_mem_inst.RAM\[38\]\[6\] _0141_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_181 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[9\].gen_latches\[5\].p_latch VGND VDPWR VDPWR
+ VGND net196 dig_ctrl_inst.latch_mem_inst.gclk\[9\] dig_ctrl_inst.latch_mem_inst.RAM\[9\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_72_48 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1922_ VDPWR VGND VDPWR VGND net133 _0582_ dig_ctrl_inst.latch_mem_inst.RAM\[32\]\[5\]
+ net50 sky130_fd_sc_hd__and3_2
X_1784_ VGND VDPWR VDPWR VGND _0444_ _0447_ _0446_ dig_ctrl_inst.latch_mem_inst.RAM\[11\]\[2\]
+ _0113_ _0445_ sky130_fd_sc_hd__a2111o_1
X_1853_ VGND VDPWR VDPWR VGND _0465_ _0515_ _0514_ sky130_fd_sc_hd__or2_1
X_2405_ VGND VDPWR VDPWR VGND _0176_ dig_ctrl_inst.spi_data_o\[5\] dig_ctrl_inst.spi_data_o\[4\]
+ _0085_ sky130_fd_sc_hd__mux2_1
X_2336_ VGND VDPWR VDPWR VGND _0958_ _0975_ _0221_ sky130_fd_sc_hd__xnor2_1
X_2198_ VDPWR VGND VDPWR VGND _0843_ _0261_ net247 _0804_ _0262_ _1039_ sky130_fd_sc_hd__o2111a_1
X_2267_ VGND VDPWR VDPWR VGND _0793_ _0909_ net161 sky130_fd_sc_hd__nor2_1
X_1218_ VGND VDPWR VDPWR VGND net248 dig_ctrl_inst.cpu_inst.instr\[6\] dig_ctrl_inst.cpu_inst.instr\[7\]
+ dig_ctrl_inst.cpu_inst.instr\[5\] _1060_ sky130_fd_sc_hd__or4b_4
Xdig_ctrl_inst.latch_mem_inst.genblk1\[5\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[5\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[5\]._gclk clknet_leaf_0_clk sky130_fd_sc_hd__dlclkp_1
Xhold31 VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.prev_state\[0\] net313 sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_data_i\[7\] net324 sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_addr\[1\] net346 sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 VGND VDPWR VDPWR VGND net19 net357 sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_addr\[5\] net335 sky130_fd_sc_hd__dlygate4sd3_1
Xhold20 VGND VDPWR VDPWR VGND dig_ctrl_inst.synchronizer_port_i_inst\[1\].pipe\[0\]
+ net302 sky130_fd_sc_hd__dlygate4sd3_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[28\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[28\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[28\]._gclk clknet_leaf_0_clk sky130_fd_sc_hd__dlclkp_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[25\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[25\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[25\]._gclk sky130_fd_sc_hd__clkbuf_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[60\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND net200 dig_ctrl_inst.latch_mem_inst.gclk\[60\] dig_ctrl_inst.latch_mem_inst.RAM\[60\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_38_276 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
XANTENNA_6 VGND VDPWR VDPWR VGND _0440_ sky130_fd_sc_hd__diode_2
X_2052_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[0\]\[7\] _0710_ _0271_
+ _0277_ sky130_fd_sc_hd__or3_1
X_2121_ VGND VDPWR VDPWR VGND net250 _1062_ net254 _0767_ sky130_fd_sc_hd__or3b_4
Xdig_ctrl_inst.latch_mem_inst.genblk1\[30\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[30\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[30\]._gclk clknet_leaf_1_clk sky130_fd_sc_hd__dlclkp_1
X_1905_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[58\]\[4\] _0158_ _0566_
+ dig_ctrl_inst.latch_mem_inst.RAM\[62\]\[4\] _0162_ sky130_fd_sc_hd__a22o_1
X_1836_ VDPWR VGND VDPWR VGND _0496_ _0494_ _0498_ _0495_ _0497_ sky130_fd_sc_hd__or4_1
X_1767_ VGND VDPWR VDPWR VGND _0430_ net101 dig_ctrl_inst.latch_mem_inst.RAM\[23\]\[2\]
+ net107 net69 sky130_fd_sc_hd__and4_1
X_1698_ VGND VDPWR VDPWR VGND _0362_ net88 dig_ctrl_inst.latch_mem_inst.RAM\[57\]\[1\]
+ net116 net41 sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_6_Right_6 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2319_ VDPWR VGND VDPWR VGND _0934_ _0959_ _0227_ sky130_fd_sc_hd__xor2_1
XFILLER_0_50_205 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xoutput21 VDPWR VGND VDPWR VGND port_ms_o[5] net21 sky130_fd_sc_hd__buf_2
Xoutput32 VDPWR VGND VDPWR VGND uo_out[7] net32 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_59_Right_59 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[53\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND net210 dig_ctrl_inst.latch_mem_inst.gclk\[53\] dig_ctrl_inst.latch_mem_inst.RAM\[53\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
X_1621_ VDPWR VGND VDPWR VGND _0280_ _0286_ _0281_ _0285_ sky130_fd_sc_hd__or3_1
X_1552_ VDPWR VGND VDPWR VGND _0218_ _1047_ _0197_ _0213_ _0025_ sky130_fd_sc_hd__a22oi_1
X_1483_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.prev_state\[0\] _0175_ dig_ctrl_inst.cpu_inst.prev_state\[1\]
+ _0174_ _1036_ _1037_ sky130_fd_sc_hd__o221ai_1
XPHY_EDGE_ROW_68_Right_68 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2104_ VGND VDPWR VDPWR VGND _0270_ _0761_ dig_ctrl_inst.cpu_inst.instr\[7\] _0034_
+ sky130_fd_sc_hd__mux2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[42\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND net223 dig_ctrl_inst.latch_mem_inst.gclk\[42\] dig_ctrl_inst.latch_mem_inst.RAM\[42\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
X_2035_ VGND VDPWR VDPWR VGND _0691_ _0694_ _0693_ dig_ctrl_inst.latch_mem_inst.RAM\[41\]\[6\]
+ _0144_ _0692_ sky130_fd_sc_hd__a2111o_1
XPHY_EDGE_ROW_77_Right_77 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1819_ VDPWR VGND VDPWR VGND net99 _0481_ dig_ctrl_inst.latch_mem_inst.RAM\[52\]\[3\]
+ net45 sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[31\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND net236 dig_ctrl_inst.latch_mem_inst.gclk\[31\] dig_ctrl_inst.latch_mem_inst.RAM\[31\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_67_113 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
Xdig_ctrl_inst.latch_mem_inst.genblk1\[5\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[5\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[5\]._gclk sky130_fd_sc_hd__clkbuf_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[57\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND net196 dig_ctrl_inst.latch_mem_inst.gclk\[57\] dig_ctrl_inst.latch_mem_inst.RAM\[57\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
Xfanout129 VGND VDPWR VDPWR VGND net130 net129 sky130_fd_sc_hd__clkbuf_2
X_2584_ VGND VDPWR VDPWR VGND net18 net173 _0098_ clknet_leaf_5_clk sky130_fd_sc_hd__dfrtp_1
Xfanout107 VGND VDPWR VDPWR VGND net108 net107 sky130_fd_sc_hd__clkbuf_2
Xfanout118 VGND VDPWR VDPWR VGND net118 net123 sky130_fd_sc_hd__clkbuf_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[46\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND net212 dig_ctrl_inst.latch_mem_inst.gclk\[46\] dig_ctrl_inst.latch_mem_inst.RAM\[46\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_1_176 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1535_ VGND VDPWR VDPWR VGND _0204_ _0185_ _0197_ _0205_ sky130_fd_sc_hd__o21ai_1
X_1604_ VGND VDPWR VDPWR VGND _0026_ _0269_ dig_ctrl_inst.cpu_inst.skip _0186_ _0266_
+ _0268_ sky130_fd_sc_hd__a32o_1
X_1466_ VDPWR VGND VDPWR VGND net265 dig_ctrl_inst.spi_data_o\[1\] dig_ctrl_inst.data_out\[1\]
+ _0164_ _1098_ sky130_fd_sc_hd__a22o_1
X_1397_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[29\] _0131_ net144
+ sky130_fd_sc_hd__and2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[35\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND net233 dig_ctrl_inst.latch_mem_inst.gclk\[35\] dig_ctrl_inst.latch_mem_inst.RAM\[35\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
X_2018_ VDPWR VGND VDPWR VGND net73 _0677_ dig_ctrl_inst.latch_mem_inst.RAM\[28\]\[6\]
+ net67 sky130_fd_sc_hd__and3_2
XFILLER_0_49_113 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[1\].gen_latches\[7\].p_latch VGND VDPWR VDPWR
+ VGND net184 dig_ctrl_inst.latch_mem_inst.gclk\[1\] dig_ctrl_inst.latch_mem_inst.RAM\[1\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[18\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[18\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[18\]._gclk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_70_119 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_51_333 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1320_ VGND VDPWR VDPWR VGND _1063_ _1158_ _1159_ _1160_ _1161_ _1162_ sky130_fd_sc_hd__o41a_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[12\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND net188 dig_ctrl_inst.latch_mem_inst.gclk\[12\] dig_ctrl_inst.latch_mem_inst.RAM\[12\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
X_1251_ VDPWR VGND VDPWR VGND net249 _1093_ net253 dig_ctrl_inst.cpu_inst.regs\[3\]\[1\]
+ sky130_fd_sc_hd__and3_2
XFILLER_0_24_85 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_24_41 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_54_193 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1518_ VGND VDPWR VDPWR VGND _0190_ dig_ctrl_inst.cpu_inst.port_o\[7\] dig_ctrl_inst.cpu_inst.regs\[0\]\[7\]
+ _0019_ sky130_fd_sc_hd__mux2_1
X_2567_ VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_receiver_inst.synchronizer_spi_cs.pipe\[0\]
+ net168 net11 clknet_leaf_4_clk sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_3 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_1449_ VDPWR VGND VDPWR VGND net84 dig_ctrl_inst.latch_mem_inst.data_we\[56\] net141
+ net37 sky130_fd_sc_hd__and3_2
X_2498_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.ip\[4\] net151 _0024_ clknet_leaf_14_clk
+ sky130_fd_sc_hd__dfrtp_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[39\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND net224 dig_ctrl_inst.latch_mem_inst.gclk\[39\] dig_ctrl_inst.latch_mem_inst.RAM\[39\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[28\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND net237 dig_ctrl_inst.latch_mem_inst.gclk\[28\] dig_ctrl_inst.latch_mem_inst.RAM\[28\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_61_17 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_51_141 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_36_160 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
Xdig_ctrl_inst.latch_mem_inst.genblk1\[35\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[35\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[35\]._gclk clknet_leaf_13_clk sky130_fd_sc_hd__dlclkp_1
XFILLER_0_36_193 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2421_ VGND VDPWR VDPWR VGND net139 dig_ctrl_inst.cpu_inst.port_o\[3\] net357 _0099_
+ sky130_fd_sc_hd__mux2_1
X_1303_ VGND VDPWR VDPWR VGND _1145_ net251 dig_ctrl_inst.cpu_inst.regs\[1\]\[5\]
+ sky130_fd_sc_hd__and2b_1
X_2283_ VDPWR VGND VDPWR VGND _1120_ _1168_ _0925_ _0877_ sky130_fd_sc_hd__a21oi_1
X_2352_ VDPWR VGND VDPWR VGND _0053_ _0990_ _0771_ _0987_ _0772_ net355 sky130_fd_sc_hd__o32a_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[16\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND net184 dig_ctrl_inst.latch_mem_inst.gclk\[16\] dig_ctrl_inst.latch_mem_inst.RAM\[16\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
X_1234_ VGND VDPWR VDPWR VGND _1076_ net249 net253 sky130_fd_sc_hd__nand2_1
X_1998_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[35\]\[6\] _0138_ _0657_
+ dig_ctrl_inst.latch_mem_inst.RAM\[53\]\[6\] _0154_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_141 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_56_17 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_72_38 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1921_ VDPWR VGND VDPWR VGND net71 _0581_ dig_ctrl_inst.latch_mem_inst.RAM\[44\]\[5\]
+ net48 sky130_fd_sc_hd__and3_2
X_1852_ VGND VDPWR VDPWR VGND _0514_ net59 dig_ctrl_inst.latch_mem_inst.RAM\[58\]\[3\]
+ _0158_ dig_ctrl_inst.latch_mem_inst.RAM\[24\]\[3\] net85 sky130_fd_sc_hd__a32o_1
X_1783_ VGND VDPWR VDPWR VGND _0446_ net76 dig_ctrl_inst.latch_mem_inst.RAM\[31\]\[2\]
+ net106 net63 sky130_fd_sc_hd__and4_1
X_2404_ VGND VDPWR VDPWR VGND _0176_ dig_ctrl_inst.spi_data_o\[4\] dig_ctrl_inst.spi_data_o\[3\]
+ _0084_ sky130_fd_sc_hd__mux2_1
X_2335_ VGND VDPWR VDPWR VGND _0974_ _0224_ _0228_ _0952_ _0973_ _0819_ sky130_fd_sc_hd__o311a_1
X_2266_ VDPWR VGND VDPWR VGND _0906_ _0908_ _0819_ _0907_ sky130_fd_sc_hd__and3_2
XFILLER_0_46_72 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_2197_ VDPWR VGND VDPWR VGND _0840_ _0842_ _0819_ _0841_ sky130_fd_sc_hd__and3_2
X_1217_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.instr\[7\] _1059_ dig_ctrl_inst.cpu_inst.instr\[6\]
+ sky130_fd_sc_hd__nor2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[61\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND net242 dig_ctrl_inst.latch_mem_inst.gclk\[61\] dig_ctrl_inst.latch_mem_inst.RAM\[61\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
Xhold32 VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.prev_state\[1\] net314 sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_receiver_inst.spi_cnt\[2\] net347
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 VGND VDPWR VDPWR VGND dig_ctrl_inst.synchronizer_mode_i_inst.pipe\[0\] net292
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 VGND VDPWR VDPWR VGND dig_ctrl_inst.synchronizer_port_i_inst\[2\].pipe\[0\]
+ net303 sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 VGND VDPWR VDPWR VGND net30 net358 sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.data\[6\] net336 sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[2\]\[1\] net325 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_225 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XANTENNA_7 VGND VDPWR VDPWR VGND _0511_ sky130_fd_sc_hd__diode_2
X_2120_ VGND VDPWR VDPWR VGND _0766_ _0764_ _0267_ _0765_ sky130_fd_sc_hd__a21o_2
X_2051_ VGND VDPWR VDPWR VGND _0270_ _0709_ dig_ctrl_inst.cpu_inst.instr\[6\] _0033_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_85 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_1904_ VDPWR VGND VDPWR VGND _0559_ _0565_ _0561_ _0564_ sky130_fd_sc_hd__or3_1
X_1835_ VGND VDPWR VDPWR VGND _0466_ _0497_ _0475_ dig_ctrl_inst.latch_mem_inst.RAM\[10\]\[3\]
+ _1190_ _0474_ sky130_fd_sc_hd__a2111o_1
X_1766_ VGND VDPWR VDPWR VGND _0429_ net103 dig_ctrl_inst.latch_mem_inst.RAM\[37\]\[2\]
+ net121 net56 sky130_fd_sc_hd__and4_1
X_1697_ VDPWR VGND VDPWR VGND net93 _0361_ dig_ctrl_inst.latch_mem_inst.RAM\[54\]\[1\]
+ net41 sky130_fd_sc_hd__and3_2
X_2318_ VGND VDPWR VDPWR VGND _0934_ _0958_ _0227_ sky130_fd_sc_hd__nor2_1
X_2249_ VGND VDPWR VDPWR VGND net163 _0892_ _0868_ sky130_fd_sc_hd__or2_1
XFILLER_0_35_203 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
Xoutput22 VDPWR VGND VDPWR VGND port_ms_o[6] net22 sky130_fd_sc_hd__buf_2
X_1482_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.prev_state\[2\] _0174_ net245
+ sky130_fd_sc_hd__xnor2_1
X_1620_ VGND VDPWR VDPWR VGND _0282_ _0285_ _0284_ dig_ctrl_inst.latch_mem_inst.RAM\[49\]\[0\]
+ _0152_ _0283_ sky130_fd_sc_hd__a2111o_1
X_1551_ VGND VDPWR VDPWR VGND _0218_ _0209_ _0185_ _0217_ dig_ctrl_inst.cpu_inst.ip\[4\]
+ dig_ctrl_inst.cpu_inst.ip\[5\] sky130_fd_sc_hd__a32o_1
X_2103_ VGND VDPWR VDPWR VGND _0761_ _0744_ _0710_ _0278_ _0760_ sky130_fd_sc_hd__o31a_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[42\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND net191 dig_ctrl_inst.latch_mem_inst.gclk\[42\] dig_ctrl_inst.latch_mem_inst.RAM\[42\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
X_2034_ VDPWR VGND VDPWR VGND net132 _0693_ dig_ctrl_inst.latch_mem_inst.RAM\[10\]\[6\]
+ net83 sky130_fd_sc_hd__and3_2
X_1818_ VDPWR VGND VDPWR VGND net73 _0480_ dig_ctrl_inst.latch_mem_inst.RAM\[28\]\[3\]
+ net63 sky130_fd_sc_hd__and3_2
XFILLER_0_4_163 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_4_141 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1749_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[15\]\[2\] _0119_ _0412_
+ dig_ctrl_inst.latch_mem_inst.RAM\[20\]\[2\] _0125_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_84 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[31\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND net203 dig_ctrl_inst.latch_mem_inst.gclk\[31\] dig_ctrl_inst.latch_mem_inst.RAM\[31\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[20\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND net223 dig_ctrl_inst.latch_mem_inst.gclk\[20\] dig_ctrl_inst.latch_mem_inst.RAM\[20\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_48_29 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[58\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND net238 dig_ctrl_inst.latch_mem_inst.gclk\[58\] dig_ctrl_inst.latch_mem_inst.RAM\[58\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_14_228 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2583_ VGND VDPWR VDPWR VGND net17 net173 _0097_ clknet_leaf_6_clk sky130_fd_sc_hd__dfrtp_1
Xfanout108 VGND VDPWR VDPWR VGND net109 net108 sky130_fd_sc_hd__clkbuf_2
X_1465_ VDPWR VGND VDPWR VGND net264 dig_ctrl_inst.spi_data_o\[0\] dig_ctrl_inst.data_out\[0\]
+ _0164_ _1080_ sky130_fd_sc_hd__a22o_1
X_2605__271 VGND VDPWR VDPWR VGND net271 _2605__271/HI sky130_fd_sc_hd__conb_1
Xfanout119 VDPWR VGND VDPWR VGND net119 net122 sky130_fd_sc_hd__buf_2
X_1534_ VDPWR VGND VDPWR VGND dig_ctrl_inst.cpu_inst.ip\[1\] _0204_ dig_ctrl_inst.cpu_inst.ip\[0\]
+ dig_ctrl_inst.cpu_inst.ip\[2\] sky130_fd_sc_hd__and3_2
X_1603_ VGND VDPWR VDPWR VGND _0269_ _0265_ net248 sky130_fd_sc_hd__nand2_1
X_2017_ VGND VDPWR VDPWR VGND _0676_ net109 dig_ctrl_inst.latch_mem_inst.RAM\[11\]\[6\]
+ net130 net90 sky130_fd_sc_hd__and4_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[42\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[42\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[42\]._gclk clknet_leaf_0_clk sky130_fd_sc_hd__dlclkp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[2\].gen_latches\[2\].p_latch VGND VDPWR VDPWR
+ VGND net220 dig_ctrl_inst.latch_mem_inst.gclk\[2\] dig_ctrl_inst.latch_mem_inst.RAM\[2\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[46\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND net179 dig_ctrl_inst.latch_mem_inst.gclk\[46\] dig_ctrl_inst.latch_mem_inst.RAM\[46\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
X_1396_ VDPWR VGND VDPWR VGND net75 _0131_ net117 net60 sky130_fd_sc_hd__and3_2
X_2612__275 VGND VDPWR VDPWR VGND net275 _2612__275/HI sky130_fd_sc_hd__conb_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[57\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[57\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[57\]._gclk sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_19_Left_97 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[35\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND net196 dig_ctrl_inst.latch_mem_inst.gclk\[35\] dig_ctrl_inst.latch_mem_inst.RAM\[35\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[24\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND net214 dig_ctrl_inst.latch_mem_inst.gclk\[24\] dig_ctrl_inst.latch_mem_inst.RAM\[24\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[13\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND net229 dig_ctrl_inst.latch_mem_inst.gclk\[13\] dig_ctrl_inst.latch_mem_inst.RAM\[13\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
X_1250_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.ip\[1\] _1073_ _1071_ _1053_
+ _1092_ sky130_fd_sc_hd__o211a_1
X_1517_ VGND VDPWR VDPWR VGND _0190_ dig_ctrl_inst.cpu_inst.port_o\[6\] net361 _0018_
+ sky130_fd_sc_hd__mux2_1
X_2566_ VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_receiver_inst.spi_mosi_sync net168
+ net299 clknet_leaf_4_clk sky130_fd_sc_hd__dfrtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[6\].gen_latches\[3\].p_latch VGND VDPWR VDPWR
+ VGND net217 dig_ctrl_inst.latch_mem_inst.gclk\[6\] dig_ctrl_inst.latch_mem_inst.RAM\[6\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
X_2497_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.ip\[3\] net152 _0023_ clknet_leaf_10_clk
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_63 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1448_ VDPWR VGND VDPWR VGND _0156_ net37 net84 sky130_fd_sc_hd__and2_1
X_1379_ VGND VDPWR VDPWR VGND net138 net104 net61 _0124_ sky130_fd_sc_hd__and3_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[39\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND net190 dig_ctrl_inst.latch_mem_inst.gclk\[39\] dig_ctrl_inst.latch_mem_inst.RAM\[39\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[28\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND net209 dig_ctrl_inst.latch_mem_inst.gclk\[28\] dig_ctrl_inst.latch_mem_inst.RAM\[28\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[17\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND net225 dig_ctrl_inst.latch_mem_inst.gclk\[17\] dig_ctrl_inst.latch_mem_inst.RAM\[17\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
X_2420_ VGND VDPWR VDPWR VGND net139 dig_ctrl_inst.cpu_inst.port_o\[2\] net18 _0098_
+ sky130_fd_sc_hd__mux2_1
Xfanout90 VDPWR VGND VDPWR VGND net90 net91 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_23_Left_101 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1233_ VGND VDPWR VDPWR VGND _1075_ _1070_ _1055_ sky130_fd_sc_hd__nand2_1
X_1302_ VDPWR VGND VDPWR VGND net251 _1144_ net255 dig_ctrl_inst.cpu_inst.regs\[3\]\[5\]
+ sky130_fd_sc_hd__and3_2
X_2282_ VDPWR VGND VDPWR VGND _1168_ _0924_ _1120_ _0877_ sky130_fd_sc_hd__and3_2
X_2351_ VGND VDPWR VDPWR VGND _0989_ _0767_ _0988_ _0990_ _0768_ sky130_fd_sc_hd__a2bb2o_1
XPHY_EDGE_ROW_32_Left_110 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1997_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[3\]\[6\] _1180_ _0656_
+ dig_ctrl_inst.latch_mem_inst.RAM\[63\]\[6\] _0163_ sky130_fd_sc_hd__a22o_1
X_2549_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[3\]\[3\] net152 _0073_
+ clknet_leaf_12_clk sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_337 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1851_ VDPWR VGND VDPWR VGND _0511_ _0509_ _0513_ _0510_ _0512_ sky130_fd_sc_hd__or4_1
X_1920_ VDPWR VGND VDPWR VGND net74 _0580_ dig_ctrl_inst.latch_mem_inst.RAM\[60\]\[5\]
+ net45 sky130_fd_sc_hd__and3_2
X_2403_ VGND VDPWR VDPWR VGND _0176_ dig_ctrl_inst.spi_data_o\[3\] dig_ctrl_inst.spi_data_o\[2\]
+ _0083_ sky130_fd_sc_hd__mux2_1
X_1782_ VGND VDPWR VDPWR VGND _0445_ net106 dig_ctrl_inst.latch_mem_inst.RAM\[19\]\[2\]
+ net136 net63 sky130_fd_sc_hd__and4_1
X_2334_ VGND VDPWR VDPWR VGND _0952_ _0228_ _0224_ _0973_ sky130_fd_sc_hd__o21ai_1
X_2196_ VDPWR VGND VDPWR VGND _1081_ _0841_ _1088_ _0263_ sky130_fd_sc_hd__or3_1
X_2265_ VGND VDPWR VDPWR VGND _0907_ _0239_ _0236_ _0889_ sky130_fd_sc_hd__a21bo_1
X_1216_ VDPWR VGND VDPWR VGND _1057_ _1058_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_320 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xhold11 VGND VDPWR VDPWR VGND dig_ctrl_inst.synchronizer_port_i_inst\[4\].pipe\[0\]
+ net293 sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 VGND VDPWR VDPWR VGND dig_ctrl_inst.stb_d net304 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[3\]\[4\] net315 sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_data_i\[0\] net337 sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[0\]\[2\] net359 sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[2\]\[0\] net326 sky130_fd_sc_hd__dlygate4sd3_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[61\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND net210 dig_ctrl_inst.latch_mem_inst.gclk\[61\] dig_ctrl_inst.latch_mem_inst.RAM\[61\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
Xhold66 VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[1\]\[3\] net348 sky130_fd_sc_hd__dlygate4sd3_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[50\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND net221 dig_ctrl_inst.latch_mem_inst.gclk\[50\] dig_ctrl_inst.latch_mem_inst.RAM\[50\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_7_Left_85 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XANTENNA_8 VGND VDPWR VDPWR VGND _1081_ sky130_fd_sc_hd__diode_2
X_2050_ VDPWR VGND VDPWR VGND _0675_ _0709_ _0708_ _0279_ dig_ctrl_inst.latch_mem_inst.RAM\[0\]\[6\]
+ sky130_fd_sc_hd__o2bb2a_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[47\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[47\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[47\]._gclk clknet_leaf_0_clk sky130_fd_sc_hd__dlclkp_1
X_1834_ VGND VDPWR VDPWR VGND _0471_ _0496_ _0487_ dig_ctrl_inst.latch_mem_inst.RAM\[15\]\[3\]
+ _0119_ _0473_ sky130_fd_sc_hd__a2111o_1
X_1903_ VGND VDPWR VDPWR VGND _0564_ _0118_ _0562_ dig_ctrl_inst.latch_mem_inst.RAM\[14\]\[4\]
+ _0563_ sky130_fd_sc_hd__a211o_1
X_1765_ VGND VDPWR VDPWR VGND _0427_ _0420_ _0428_ _0406_ _0413_ sky130_fd_sc_hd__nor4_1
XFILLER_0_32_75 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_1696_ VGND VDPWR VDPWR VGND _0360_ net103 dig_ctrl_inst.latch_mem_inst.RAM\[55\]\[1\]
+ net105 net41 sky130_fd_sc_hd__and4_1
XFILLER_0_32_3 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_2317_ VGND VDPWR VDPWR VGND _1114_ _0956_ _0859_ net162 _0957_ sky130_fd_sc_hd__o211a_1
X_2248_ VDPWR VGND VDPWR VGND _0889_ _0891_ _0819_ _0890_ sky130_fd_sc_hd__and3_2
X_2179_ VDPWR VGND VDPWR VGND dig_ctrl_inst.cpu_inst.data\[2\] dig_ctrl_inst.cpu_inst.data\[0\]
+ dig_ctrl_inst.cpu_inst.data\[3\] _0825_ _0823_ sky130_fd_sc_hd__or4b_1
Xoutput23 VDPWR VGND VDPWR VGND port_ms_o[7] net23 sky130_fd_sc_hd__buf_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[54\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND net211 dig_ctrl_inst.latch_mem_inst.gclk\[54\] dig_ctrl_inst.latch_mem_inst.RAM\[54\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_34_270 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_109 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1481_ VDPWR VGND VDPWR VGND _1036_ dig_ctrl_inst.cpu_inst.prev_state\[0\] _0173_
+ _1037_ dig_ctrl_inst.cpu_inst.prev_state\[1\] sky130_fd_sc_hd__a22o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[43\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND net233 dig_ctrl_inst.latch_mem_inst.gclk\[43\] dig_ctrl_inst.latch_mem_inst.RAM\[43\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[21\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[21\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[21\]._gclk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_337 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1550_ VDPWR VGND VDPWR VGND _0216_ _0217_ sky130_fd_sc_hd__inv_2
X_2102_ VDPWR VGND VDPWR VGND _0755_ _0747_ _0760_ _0750_ _0759_ sky130_fd_sc_hd__or4_1
X_2033_ VDPWR VGND VDPWR VGND net111 _0692_ dig_ctrl_inst.latch_mem_inst.RAM\[34\]\[6\]
+ net52 sky130_fd_sc_hd__and3_2
X_1817_ VGND VDPWR VDPWR VGND _0479_ net107 dig_ctrl_inst.latch_mem_inst.RAM\[11\]\[3\]
+ net131 net91 sky130_fd_sc_hd__and4_1
X_1748_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[1\]\[2\] _1175_ _0411_
+ dig_ctrl_inst.latch_mem_inst.RAM\[2\]\[2\] _1178_ sky130_fd_sc_hd__a22o_1
X_1679_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[2\]\[1\] _1178_ _0343_
+ dig_ctrl_inst.latch_mem_inst.RAM\[60\]\[1\] _0160_ sky130_fd_sc_hd__a22o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[20\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND net192 dig_ctrl_inst.latch_mem_inst.gclk\[20\] dig_ctrl_inst.latch_mem_inst.RAM\[20\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[58\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND net205 dig_ctrl_inst.latch_mem_inst.gclk\[58\] dig_ctrl_inst.latch_mem_inst.RAM\[58\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
X_2582_ VGND VDPWR VDPWR VGND net16 net173 _0096_ clknet_leaf_6_clk sky130_fd_sc_hd__dfrtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[47\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND net223 dig_ctrl_inst.latch_mem_inst.gclk\[47\] dig_ctrl_inst.latch_mem_inst.RAM\[47\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
X_1602_ VDPWR VGND VDPWR VGND dig_ctrl_inst.cpu_inst.instr\[7\] _0268_ dig_ctrl_inst.cpu_inst.instr\[6\]
+ _0189_ sky130_fd_sc_hd__and3_2
Xfanout109 VDPWR VGND VDPWR VGND net109 net110 sky130_fd_sc_hd__buf_2
X_1464_ VDPWR VGND VDPWR VGND _1041_ _0164_ net167 sky130_fd_sc_hd__and2_2
X_1395_ VDPWR VGND VDPWR VGND net73 dig_ctrl_inst.latch_mem_inst.data_we\[28\] net145
+ net67 sky130_fd_sc_hd__and3_2
X_1533_ VGND VDPWR VDPWR VGND _0197_ _0203_ dig_ctrl_inst.cpu_inst.ip\[1\] _0021_
+ sky130_fd_sc_hd__mux2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[36\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND net238 dig_ctrl_inst.latch_mem_inst.gclk\[36\] dig_ctrl_inst.latch_mem_inst.RAM\[36\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_49_137 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[2\].gen_latches\[6\].p_latch VGND VDPWR VDPWR
+ VGND net186 dig_ctrl_inst.latch_mem_inst.gclk\[2\] dig_ctrl_inst.latch_mem_inst.RAM\[2\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
X_2016_ VGND VDPWR VDPWR VGND _0674_ _0667_ _0675_ _0655_ _0660_ sky130_fd_sc_hd__nor4_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[24\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND net179 dig_ctrl_inst.latch_mem_inst.gclk\[24\] dig_ctrl_inst.latch_mem_inst.RAM\[24\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[13\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND net195 dig_ctrl_inst.latch_mem_inst.gclk\[13\] dig_ctrl_inst.latch_mem_inst.RAM\[13\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_20_Left_98 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_12_clk VGND VDPWR VDPWR VGND clknet_leaf_12_clk clknet_1_0__leaf_clk
+ sky130_fd_sc_hd__clkbuf_8
X_1516_ VGND VDPWR VDPWR VGND _0190_ dig_ctrl_inst.cpu_inst.port_o\[5\] net343 _0017_
+ sky130_fd_sc_hd__mux2_1
X_2565_ VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_receiver_inst.synchronizer_spi_mosi.pipe\[0\]
+ net168 net12 clknet_leaf_4_clk sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_64 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_1447_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[55\] _0155_ net148
+ sky130_fd_sc_hd__and2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[6\].gen_latches\[7\].p_latch VGND VDPWR VDPWR
+ VGND net180 dig_ctrl_inst.latch_mem_inst.gclk\[6\] dig_ctrl_inst.latch_mem_inst.RAM\[6\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[1\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[1\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[1\]._gclk sky130_fd_sc_hd__clkbuf_4
X_2496_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.ip\[2\] net153 _0022_ clknet_leaf_10_clk
+ sky130_fd_sc_hd__dfrtp_2
X_1378_ VDPWR VGND VDPWR VGND net111 dig_ctrl_inst.latch_mem_inst.data_we\[18\] net141
+ net61 sky130_fd_sc_hd__and3_2
XFILLER_0_5_292 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
Xfanout91 VDPWR VGND VDPWR VGND net91 net92 sky130_fd_sc_hd__buf_2
Xfanout80 VGND VDPWR VDPWR VGND _0114_ net80 sky130_fd_sc_hd__clkbuf_2
Xdig_ctrl_inst.latch_mem_inst.genblk1\[14\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[14\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[14\]._gclk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_36_151 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_28_118 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
Xdig_ctrl_inst.latch_mem_inst.gen_words\[17\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND net190 dig_ctrl_inst.latch_mem_inst.gclk\[17\] dig_ctrl_inst.latch_mem_inst.RAM\[17\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_36_173 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_1301_ VGND VDPWR VDPWR VGND net255 net251 _1143_ dig_ctrl_inst.cpu_inst.regs\[2\]\[5\]
+ sky130_fd_sc_hd__and3b_1
X_2350_ VDPWR VGND VDPWR VGND dig_ctrl_inst.spi_data_o\[7\] _0183_ _0989_ dig_ctrl_inst.synchronizer_port_i_inst\[7\].out
+ _0824_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_1_clk VGND VDPWR VDPWR VGND clknet_leaf_1_clk clknet_1_1__leaf_clk sky130_fd_sc_hd__clkbuf_8
X_2281_ VDPWR VGND VDPWR VGND _0912_ _1114_ _0922_ _0923_ sky130_fd_sc_hd__a21o_1
X_1232_ VGND VDPWR VDPWR VGND _1074_ _1070_ _1072_ _1054_ _1040_ sky130_fd_sc_hd__a211o_1
XFILLER_0_19_107 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_51_52 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1996_ VDPWR VGND VDPWR VGND _0649_ _0655_ _0650_ _0654_ sky130_fd_sc_hd__or3_1
XFILLER_0_15_324 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_3 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2548_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[3\]\[2\] net154 _0072_
+ clknet_leaf_12_clk sky130_fd_sc_hd__dfrtp_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[54\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[54\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[54\]._gclk clknet_leaf_16_clk sky130_fd_sc_hd__dlclkp_1
X_2479_ VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_data_i\[1\] net173 _0005_ clknet_leaf_5_clk
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_165 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xclkload0 VGND VDPWR VDPWR VGND clknet_1_0__leaf_clk clkload0/Y sky130_fd_sc_hd__inv_8
XFILLER_0_33_187 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_305 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1850_ VGND VDPWR VDPWR VGND _0478_ _0512_ _0493_ dig_ctrl_inst.latch_mem_inst.RAM\[7\]\[3\]
+ _1184_ _0491_ sky130_fd_sc_hd__a2111o_1
X_1781_ VDPWR VGND VDPWR VGND net86 _0444_ dig_ctrl_inst.latch_mem_inst.RAM\[40\]\[2\]
+ net53 sky130_fd_sc_hd__and3_2
X_2402_ VGND VDPWR VDPWR VGND _0176_ dig_ctrl_inst.spi_data_o\[2\] dig_ctrl_inst.spi_data_o\[1\]
+ _0082_ sky130_fd_sc_hd__mux2_1
X_2333_ VDPWR VGND VDPWR VGND _0052_ _0972_ _0771_ _0967_ _0772_ net354 sky130_fd_sc_hd__o32a_1
XFILLER_0_46_41 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2264_ VGND VDPWR VDPWR VGND _0236_ _0889_ _0906_ _0238_ sky130_fd_sc_hd__or3b_1
X_2195_ VGND VDPWR VDPWR VGND _0840_ _0263_ _0259_ sky130_fd_sc_hd__nand2_1
X_1215_ VGND VDPWR VDPWR VGND net249 _1057_ net253 sky130_fd_sc_hd__nand2b_2
XFILLER_0_62_216 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1979_ VGND VDPWR VDPWR VGND _0581_ _0639_ _0622_ dig_ctrl_inst.latch_mem_inst.RAM\[10\]\[5\]
+ _1190_ _0602_ sky130_fd_sc_hd__a2111o_1
Xhold12 VGND VDPWR VDPWR VGND dig_ctrl_inst.synchronizer_port_ms_i_inst.pipe\[0\]
+ net294 sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[2\]\[6\] net338 sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 VGND VDPWR VDPWR VGND net21 net327 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_receiver_inst.spi_sclk_sync net305
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[1\]\[5\] net316 sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[0\]\[3\] net349 sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 VGND VDPWR VDPWR VGND net29 net360 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_51_Left_129 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_60_Left_138 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[50\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND net194 dig_ctrl_inst.latch_mem_inst.gclk\[50\] dig_ctrl_inst.latch_mem_inst.RAM\[50\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
XANTENNA_9 VGND VDPWR VDPWR VGND _1173_ sky130_fd_sc_hd__diode_2
X_1902_ VDPWR VGND VDPWR VGND _0563_ _0272_ dig_ctrl_inst.latch_mem_inst.RAM\[10\]\[4\]
+ dig_ctrl_inst.latch_mem_inst.RAM\[5\]\[4\] _1190_ _0539_ sky130_fd_sc_hd__a221o_1
X_1833_ VGND VDPWR VDPWR VGND _0468_ _0495_ _0488_ dig_ctrl_inst.latch_mem_inst.RAM\[1\]\[3\]
+ _1175_ _0483_ sky130_fd_sc_hd__a2111o_1
X_1764_ VDPWR VGND VDPWR VGND _0424_ _0427_ _0425_ _0426_ sky130_fd_sc_hd__or3_1
X_1695_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[11\]\[1\] _0113_ _0359_
+ dig_ctrl_inst.latch_mem_inst.RAM\[27\]\[1\] _0130_ sky130_fd_sc_hd__a22o_1
X_2316_ VDPWR VGND VDPWR VGND _0954_ _0862_ _0956_ _0909_ _0955_ sky130_fd_sc_hd__or4_1
XFILLER_0_12_179 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2247_ VGND VDPWR VDPWR VGND _0890_ _0241_ _0872_ _0244_ sky130_fd_sc_hd__nand3_1
X_2178_ VGND VDPWR VDPWR VGND _0823_ _0180_ dig_ctrl_inst.cpu_inst.data\[0\] _0824_
+ sky130_fd_sc_hd__nor3b_4
Xoutput24 VDPWR VGND VDPWR VGND uio_out[2] net24 sky130_fd_sc_hd__buf_2
Xdig_ctrl_inst.latch_mem_inst.genblk1\[60\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[60\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[60\]._gclk sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_19_Right_19 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[54\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND net184 dig_ctrl_inst.latch_mem_inst.gclk\[54\] dig_ctrl_inst.latch_mem_inst.RAM\[54\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_1_305 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1480_ VDPWR VGND VDPWR VGND net266 dig_ctrl_inst.spi_data_o\[7\] dig_ctrl_inst.data_out\[7\]
+ _0172_ _0164_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_10 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_28_Right_28 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[43\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND net201 dig_ctrl_inst.latch_mem_inst.gclk\[43\] dig_ctrl_inst.latch_mem_inst.RAM\[43\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
X_2101_ VDPWR VGND VDPWR VGND _0757_ _0723_ _0759_ _0756_ _0758_ sky130_fd_sc_hd__or4_1
X_2032_ VGND VDPWR VDPWR VGND _0691_ net76 dig_ctrl_inst.latch_mem_inst.RAM\[31\]\[6\]
+ net105 net62 sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_37_Right_37 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[32\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND net211 dig_ctrl_inst.latch_mem_inst.gclk\[32\] dig_ctrl_inst.latch_mem_inst.RAM\[32\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_46_Right_46 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1816_ VGND VDPWR VDPWR VGND _0478_ net107 dig_ctrl_inst.latch_mem_inst.RAM\[51\]\[3\]
+ net136 net47 sky130_fd_sc_hd__and4_1
X_1678_ VGND VDPWR VDPWR VGND _0342_ net49 dig_ctrl_inst.latch_mem_inst.RAM\[41\]\[1\]
+ _0144_ dig_ctrl_inst.latch_mem_inst.RAM\[44\]\[1\] net71 sky130_fd_sc_hd__a32o_1
XFILLER_0_32_219 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1747_ VGND VDPWR VDPWR VGND _0407_ _0410_ _0409_ dig_ctrl_inst.latch_mem_inst.RAM\[43\]\[2\]
+ _0146_ _0408_ sky130_fd_sc_hd__a2111o_1
XPHY_EDGE_ROW_55_Right_55 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[21\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND net232 dig_ctrl_inst.latch_mem_inst.gclk\[21\] dig_ctrl_inst.latch_mem_inst.RAM\[21\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_64_Right_64 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_16_282 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_73_Right_73 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2581_ VGND VDPWR VDPWR VGND net32 net172 _0095_ clknet_leaf_6_clk sky130_fd_sc_hd__dfrtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[47\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND net191 dig_ctrl_inst.latch_mem_inst.gclk\[47\] dig_ctrl_inst.latch_mem_inst.RAM\[47\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[3\].gen_latches\[1\].p_latch VGND VDPWR VDPWR
+ VGND net232 dig_ctrl_inst.latch_mem_inst.gclk\[3\] dig_ctrl_inst.latch_mem_inst.RAM\[3\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
X_1532_ VDPWR VGND VDPWR VGND _0185_ _0201_ _0203_ _0200_ _0202_ sky130_fd_sc_hd__a22o_1
X_1601_ VGND VDPWR VDPWR VGND _0267_ dig_ctrl_inst.cpu_inst.instr\[7\] dig_ctrl_inst.cpu_inst.instr\[6\]
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_42 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.genblk1\[59\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[59\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[59\]._gclk clknet_leaf_2_clk sky130_fd_sc_hd__dlclkp_1
X_1394_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[27\] _0130_ net146
+ sky130_fd_sc_hd__and2_1
X_1463_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[63\] _0163_ net144
+ sky130_fd_sc_hd__and2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[36\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND net209 dig_ctrl_inst.latch_mem_inst.gclk\[36\] dig_ctrl_inst.latch_mem_inst.RAM\[36\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
X_2015_ VDPWR VGND VDPWR VGND _0668_ _0674_ _0669_ _0673_ sky130_fd_sc_hd__or3_1
XFILLER_0_9_246 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
Xdig_ctrl_inst.latch_mem_inst.gen_words\[25\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND net219 dig_ctrl_inst.latch_mem_inst.gclk\[25\] dig_ctrl_inst.latch_mem_inst.RAM\[25\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_input_latches\[2\].n_latch VGND VDPWR VDPWR VGND
+ dig_ctrl_inst.data_out\[2\] clknet_leaf_9_clk dig_ctrl_inst.latch_mem_inst.wdata\[2\]
+ sky130_fd_sc_hd__dlxtn_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[61\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[61\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[61\]._gclk clknet_leaf_2_clk sky130_fd_sc_hd__dlclkp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[14\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND net240 dig_ctrl_inst.latch_mem_inst.gclk\[14\] dig_ctrl_inst.latch_mem_inst.RAM\[14\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[7\].gen_latches\[2\].p_latch VGND VDPWR VDPWR
+ VGND net226 dig_ctrl_inst.latch_mem_inst.gclk\[7\] dig_ctrl_inst.latch_mem_inst.RAM\[7\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_27_333 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1515_ VGND VDPWR VDPWR VGND _0190_ dig_ctrl_inst.cpu_inst.port_o\[4\] net341 _0016_
+ sky130_fd_sc_hd__mux2_1
X_2564_ VDPWR VGND VDPWR VGND dig_ctrl_inst.spi_receiver_inst.spi_sclk_delayed clknet_leaf_4_clk
+ net305 sky130_fd_sc_hd__dfxtp_1
X_2495_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.ip\[1\] net153 _0021_ clknet_leaf_14_clk
+ sky130_fd_sc_hd__dfrtp_1
X_1446_ VDPWR VGND VDPWR VGND net102 _0155_ net106 net43 sky130_fd_sc_hd__and3_2
X_1377_ VDPWR VGND VDPWR VGND _0123_ net63 net113 sky130_fd_sc_hd__and2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[29\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND net213 dig_ctrl_inst.latch_mem_inst.gclk\[29\] dig_ctrl_inst.latch_mem_inst.RAM\[29\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[53\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[53\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[53\]._gclk sky130_fd_sc_hd__clkbuf_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[18\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND net231 dig_ctrl_inst.latch_mem_inst.gclk\[18\] dig_ctrl_inst.latch_mem_inst.RAM\[18\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
Xfanout70 VGND VDPWR VDPWR VGND _0120_ net70 sky130_fd_sc_hd__clkbuf_2
Xfanout92 VGND VDPWR VDPWR VGND _1185_ net92 sky130_fd_sc_hd__clkbuf_2
Xfanout81 VDPWR VGND VDPWR VGND net81 net83 sky130_fd_sc_hd__buf_2
XFILLER_0_36_141 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_36_185 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_10_24 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2280_ VGND VDPWR VDPWR VGND _0921_ _0920_ _0922_ _0908_ sky130_fd_sc_hd__or3b_1
X_1300_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.ip\[5\] _1073_ _1071_ _1053_
+ _1142_ sky130_fd_sc_hd__o211a_1
X_1231_ VGND VDPWR VDPWR VGND _1073_ _1054_ _1056_ sky130_fd_sc_hd__nand2_2
X_1995_ VGND VDPWR VDPWR VGND _0651_ _0654_ _0653_ dig_ctrl_inst.latch_mem_inst.RAM\[59\]\[6\]
+ _0159_ _0652_ sky130_fd_sc_hd__a2111o_1
X_2478_ VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_data_i\[0\] net173 _0004_ clknet_leaf_6_clk
+ sky130_fd_sc_hd__dfrtp_1
X_1429_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[45\] _0147_ net146
+ sky130_fd_sc_hd__and2_1
X_2547_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[3\]\[1\] net155 _0071_
+ clknet_leaf_12_clk sky130_fd_sc_hd__dfrtp_1
Xclkload1 VGND VDPWR VDPWR VGND clkload1/Y clknet_leaf_10_clk sky130_fd_sc_hd__inv_16
XFILLER_0_33_144 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_33_199 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
Xfanout260 VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.arg0\[1\] net260 sky130_fd_sc_hd__clkbuf_2
X_1780_ VGND VDPWR VDPWR VGND _0442_ _0440_ _0443_ _0432_ _0436_ sky130_fd_sc_hd__nor4_1
XFILLER_0_21_23 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_24_177 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_2401_ VGND VDPWR VDPWR VGND _0176_ dig_ctrl_inst.spi_data_o\[1\] dig_ctrl_inst.spi_data_o\[0\]
+ _0081_ sky130_fd_sc_hd__mux2_1
X_2332_ VGND VDPWR VDPWR VGND _0971_ _0767_ _0970_ _0972_ _0768_ sky130_fd_sc_hd__a2bb2o_1
X_2194_ VGND VDPWR VDPWR VGND _0839_ _0797_ _0836_ _0838_ _0833_ _1114_ sky130_fd_sc_hd__o311a_1
X_2263_ VDPWR VGND VDPWR VGND _0049_ _0905_ _0771_ _0902_ _0772_ net349 sky130_fd_sc_hd__o32a_1
X_1214_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.cpu_state\[0\] dig_ctrl_inst.cpu_inst.cpu_state\[1\]
+ _1056_ net245 sky130_fd_sc_hd__or3b_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[62\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND net213 dig_ctrl_inst.latch_mem_inst.gclk\[62\] dig_ctrl_inst.latch_mem_inst.RAM\[62\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
X_1978_ VGND VDPWR VDPWR VGND _0616_ _0638_ _0624_ dig_ctrl_inst.latch_mem_inst.RAM\[15\]\[5\]
+ _0119_ _0619_ sky130_fd_sc_hd__a2111o_1
Xhold68 VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_data_o\[7\] net350 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[0\]\[6\] net361 sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 VGND VDPWR VDPWR VGND net22 net328 sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_data_i\[4\] net317 sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 VGND VDPWR VDPWR VGND dig_ctrl_inst.mode_sync net306 sky130_fd_sc_hd__dlygate4sd3_1
Xhold13 VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_receiver_inst.synchronizer_spi_cs.pipe\[0\]
+ net295 sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[2\]\[3\] net339 sky130_fd_sc_hd__dlygate4sd3_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[51\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND net234 dig_ctrl_inst.latch_mem_inst.gclk\[51\] dig_ctrl_inst.latch_mem_inst.RAM\[51\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_46_280 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_21_136 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1832_ VDPWR VGND VDPWR VGND _0494_ _0142_ dig_ctrl_inst.latch_mem_inst.RAM\[38\]\[3\]
+ dig_ctrl_inst.latch_mem_inst.RAM\[39\]\[3\] _0141_ _0481_ sky130_fd_sc_hd__a221o_1
X_1901_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[29\]\[4\] _0131_ _0562_
+ dig_ctrl_inst.latch_mem_inst.RAM\[33\]\[4\] _0136_ sky130_fd_sc_hd__a22o_1
X_1694_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[29\]\[1\] _0131_ _0358_
+ dig_ctrl_inst.latch_mem_inst.RAM\[58\]\[1\] _0158_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_336 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
X_1763_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[48\]\[2\] _0151_ _0426_
+ dig_ctrl_inst.latch_mem_inst.RAM\[63\]\[2\] _0163_ sky130_fd_sc_hd__a22o_1
X_2246_ VDPWR VGND VDPWR VGND _0872_ _0244_ _0241_ _0889_ sky130_fd_sc_hd__a21o_1
X_2315_ VGND VDPWR VDPWR VGND _0794_ _0784_ _0779_ _1081_ _0955_ sky130_fd_sc_hd__o211a_1
XFILLER_0_73_51 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2177_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.data\[1\] _0823_ _0181_ sky130_fd_sc_hd__or2_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[46\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[46\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[46\]._gclk sky130_fd_sc_hd__clkbuf_4
Xoutput25 VDPWR VGND VDPWR VGND uo_out[0] net25 sky130_fd_sc_hd__buf_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[55\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND net220 dig_ctrl_inst.latch_mem_inst.gclk\[55\] dig_ctrl_inst.latch_mem_inst.RAM\[55\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[44\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND net242 dig_ctrl_inst.latch_mem_inst.gclk\[44\] dig_ctrl_inst.latch_mem_inst.RAM\[44\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
X_2100_ VGND VDPWR VDPWR VGND _0758_ net63 dig_ctrl_inst.latch_mem_inst.RAM\[18\]\[7\]
+ _0123_ dig_ctrl_inst.latch_mem_inst.RAM\[28\]\[7\] net72 sky130_fd_sc_hd__a32o_1
X_2031_ VGND VDPWR VDPWR VGND _0689_ _0685_ _0690_ _0679_ _0683_ sky130_fd_sc_hd__nor4_1
X_1815_ VGND VDPWR VDPWR VGND _0477_ net76 dig_ctrl_inst.latch_mem_inst.RAM\[62\]\[3\]
+ net114 net41 sky130_fd_sc_hd__and4_1
XFILLER_0_32_209 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_4_100 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_68_62 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1677_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[9\]\[1\] _1188_ _0341_
+ dig_ctrl_inst.latch_mem_inst.RAM\[10\]\[1\] _1190_ sky130_fd_sc_hd__a22o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[32\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND net179 dig_ctrl_inst.latch_mem_inst.gclk\[32\] dig_ctrl_inst.latch_mem_inst.RAM\[32\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
X_1746_ VDPWR VGND VDPWR VGND net111 _0409_ dig_ctrl_inst.latch_mem_inst.RAM\[50\]\[2\]
+ net40 sky130_fd_sc_hd__and3_2
X_2229_ VGND VDPWR VDPWR VGND _0873_ _0872_ _0819_ sky130_fd_sc_hd__nand2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[21\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND net202 dig_ctrl_inst.latch_mem_inst.gclk\[21\] dig_ctrl_inst.latch_mem_inst.RAM\[21\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_16_294 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
Xdig_ctrl_inst.latch_mem_inst.gen_words\[59\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND net217 dig_ctrl_inst.latch_mem_inst.gclk\[59\] dig_ctrl_inst.latch_mem_inst.RAM\[59\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[10\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND net211 dig_ctrl_inst.latch_mem_inst.gclk\[10\] dig_ctrl_inst.latch_mem_inst.RAM\[10\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_7_3 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
Xdig_ctrl_inst.latch_mem_inst.gen_words\[48\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND net235 dig_ctrl_inst.latch_mem_inst.gclk\[48\] dig_ctrl_inst.latch_mem_inst.RAM\[48\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_13_57 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1462_ VDPWR VGND VDPWR VGND net75 _0163_ net104 net39 sky130_fd_sc_hd__and3_2
X_2580_ VGND VDPWR VDPWR VGND net31 net172 _0094_ clknet_leaf_6_clk sky130_fd_sc_hd__dfrtp_1
X_1600_ VGND VDPWR VDPWR VGND net248 _0266_ _0265_ sky130_fd_sc_hd__or2_1
X_1531_ VGND VDPWR VDPWR VGND _0202_ dig_ctrl_inst.cpu_inst.ip\[0\] _0186_ dig_ctrl_inst.cpu_inst.ip\[1\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_38_54 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[3\].gen_latches\[5\].p_latch VGND VDPWR VDPWR
+ VGND net201 dig_ctrl_inst.latch_mem_inst.gclk\[3\] dig_ctrl_inst.latch_mem_inst.RAM\[3\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
X_1393_ VDPWR VGND VDPWR VGND net90 _0130_ net109 net67 sky130_fd_sc_hd__and3_2
XFILLER_0_9_258 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
X_2014_ VGND VDPWR VDPWR VGND _0670_ _0673_ _0672_ dig_ctrl_inst.latch_mem_inst.RAM\[19\]\[6\]
+ _0124_ _0671_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_13_220 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1729_ VDPWR VGND VDPWR VGND net94 _0393_ dig_ctrl_inst.latch_mem_inst.RAM\[22\]\[1\]
+ net65 sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_input_latches\[6\].n_latch VGND VDPWR VDPWR VGND
+ dig_ctrl_inst.data_out\[6\] clknet_leaf_9_clk dig_ctrl_inst.latch_mem_inst.wdata\[6\]
+ sky130_fd_sc_hd__dlxtn_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[25\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND net186 dig_ctrl_inst.latch_mem_inst.gclk\[25\] dig_ctrl_inst.latch_mem_inst.RAM\[25\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[14\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND net203 dig_ctrl_inst.latch_mem_inst.gclk\[14\] dig_ctrl_inst.latch_mem_inst.RAM\[14\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_51_337 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_39_161 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1514_ VGND VDPWR VDPWR VGND _0190_ dig_ctrl_inst.cpu_inst.port_o\[3\] net349 _0015_
+ sky130_fd_sc_hd__mux2_1
X_2563_ VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_data_o\[7\] net171 net351 clknet_leaf_3_clk
+ sky130_fd_sc_hd__dfrtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[7\].gen_latches\[6\].p_latch VGND VDPWR VDPWR
+ VGND net193 dig_ctrl_inst.latch_mem_inst.gclk\[7\] dig_ctrl_inst.latch_mem_inst.RAM\[7\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_49_31 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2494_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.ip\[0\] net153 _0020_ clknet_leaf_14_clk
+ sky130_fd_sc_hd__dfrtp_1
X_1445_ VDPWR VGND VDPWR VGND net93 dig_ctrl_inst.latch_mem_inst.data_we\[54\] net141
+ net37 sky130_fd_sc_hd__and3_2
X_1376_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[17\] _0122_ net147
+ sky130_fd_sc_hd__and2_1
XFILLER_0_65_41 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
Xdig_ctrl_inst.latch_mem_inst.genblk1\[39\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[39\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[39\]._gclk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_37_109 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_45_164 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[29\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND net178 dig_ctrl_inst.latch_mem_inst.gclk\[29\] dig_ctrl_inst.latch_mem_inst.RAM\[29\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[18\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND net195 dig_ctrl_inst.latch_mem_inst.gclk\[18\] dig_ctrl_inst.latch_mem_inst.RAM\[18\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
Xfanout82 VGND VDPWR VDPWR VGND net83 net82 sky130_fd_sc_hd__clkbuf_2
Xfanout93 VDPWR VGND VDPWR VGND net93 net96 sky130_fd_sc_hd__buf_2
Xfanout60 VGND VDPWR VDPWR VGND net61 net60 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_36_197 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xfanout71 VDPWR VGND VDPWR VGND net71 _0115_ sky130_fd_sc_hd__buf_2
X_1230_ VGND VDPWR VDPWR VGND _1055_ _1072_ _1053_ sky130_fd_sc_hd__nor2_1
X_1994_ VDPWR VGND VDPWR VGND net113 _0653_ dig_ctrl_inst.latch_mem_inst.RAM\[50\]\[6\]
+ net46 sky130_fd_sc_hd__and3_2
X_2615_ VDPWR VGND VDPWR VGND uio_out[7] net278 sky130_fd_sc_hd__buf_2
XFILLER_0_15_337 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2546_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[3\]\[0\] net156 _0070_
+ clknet_leaf_8_clk sky130_fd_sc_hd__dfrtp_1
X_2477_ VGND VDPWR VDPWR VGND dig_ctrl_inst.port_ms_sync_i net175 net294 clknet_leaf_8_clk
+ sky130_fd_sc_hd__dfrtp_1
X_1428_ VDPWR VGND VDPWR VGND net79 _0147_ net120 net55 sky130_fd_sc_hd__and3_2
X_1359_ VDPWR VGND VDPWR VGND net142 dig_ctrl_inst.latch_mem_inst.data_we\[10\] net126
+ net83 sky130_fd_sc_hd__and3_2
Xclkload2 VGND VDPWR VDPWR VGND clkload2/Y clknet_leaf_11_clk sky130_fd_sc_hd__inv_16
Xfanout250 VDPWR VGND VDPWR VGND net250 net252 sky130_fd_sc_hd__buf_2
Xfanout261 VGND VDPWR VDPWR VGND net263 net261 sky130_fd_sc_hd__clkbuf_2
X_2400_ VGND VDPWR VDPWR VGND _0176_ dig_ctrl_inst.spi_data_o\[0\] net307 _0080_ sky130_fd_sc_hd__mux2_1
X_1213_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.cpu_state\[1\] _1055_ dig_ctrl_inst.cpu_inst.cpu_state\[0\]
+ net245 sky130_fd_sc_hd__nor3b_2
X_2331_ VDPWR VGND VDPWR VGND dig_ctrl_inst.spi_data_o\[6\] _0183_ _0971_ dig_ctrl_inst.synchronizer_port_i_inst\[6\].out
+ _0824_ sky130_fd_sc_hd__a22o_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[10\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[10\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[10\]._gclk sky130_fd_sc_hd__clkbuf_4
X_2262_ VGND VDPWR VDPWR VGND _0904_ _0767_ _0903_ _0905_ _0768_ sky130_fd_sc_hd__a2bb2o_1
X_2193_ VGND VDPWR VDPWR VGND _0834_ _0837_ _0838_ _0782_ _0776_ sky130_fd_sc_hd__o22ai_1
X_1977_ VGND VDPWR VDPWR VGND _0615_ _0637_ _0623_ dig_ctrl_inst.latch_mem_inst.RAM\[62\]\[5\]
+ _0162_ _0621_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_30_126 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_2529_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[1\]\[1\] net152 _0055_
+ clknet_leaf_12_clk sky130_fd_sc_hd__dfrtp_1
Xhold14 VGND VDPWR VDPWR VGND dig_ctrl_inst.synchronizer_port_i_inst\[7\].pipe\[0\]
+ net296 sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_receiver_inst.spi_mosi_sync net307
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 VGND VDPWR VDPWR VGND _0087_ net351 sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[1\]\[4\] net340 sky130_fd_sc_hd__dlygate4sd3_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[62\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND net178 dig_ctrl_inst.latch_mem_inst.gclk\[62\] dig_ctrl_inst.latch_mem_inst.RAM\[62\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
Xhold36 VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[3\]\[1\] net318 sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.data\[7\] net329 sky130_fd_sc_hd__dlygate4sd3_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[51\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND net200 dig_ctrl_inst.latch_mem_inst.gclk\[51\] dig_ctrl_inst.latch_mem_inst.RAM\[51\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[40\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND net213 dig_ctrl_inst.latch_mem_inst.gclk\[40\] dig_ctrl_inst.latch_mem_inst.RAM\[40\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_44_218 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
X_1831_ VDPWR VGND VDPWR VGND net99 _0493_ dig_ctrl_inst.latch_mem_inst.RAM\[20\]\[3\]
+ net69 sky130_fd_sc_hd__and3_2
X_1900_ VDPWR VGND VDPWR VGND _0561_ _0144_ dig_ctrl_inst.latch_mem_inst.RAM\[9\]\[4\]
+ dig_ctrl_inst.latch_mem_inst.RAM\[41\]\[4\] _1188_ _0560_ sky130_fd_sc_hd__a221o_1
X_2608__272 VGND VDPWR VDPWR VGND net272 _2608__272/HI sky130_fd_sc_hd__conb_1
X_1693_ VDPWR VGND VDPWR VGND _0354_ _0357_ _0355_ _0356_ sky130_fd_sc_hd__or3_1
X_1762_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[14\]\[2\] _0118_ _0425_
+ dig_ctrl_inst.latch_mem_inst.RAM\[25\]\[2\] _0129_ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_53 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2245_ VGND VDPWR VDPWR VGND _1114_ _0886_ _0887_ net162 _0888_ sky130_fd_sc_hd__o211a_1
X_2176_ VDPWR VGND VDPWR VGND _0811_ _0822_ _0803_ _0821_ sky130_fd_sc_hd__and3_2
X_2314_ VGND VDPWR VDPWR VGND _0910_ _0954_ _0857_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_142 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xoutput26 VDPWR VGND VDPWR VGND uo_out[1] net26 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_1_Right_1 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xoutput15 VGND VDPWR VDPWR VGND clk_o net15 sky130_fd_sc_hd__clkbuf_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[55\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND net190 dig_ctrl_inst.latch_mem_inst.gclk\[55\] dig_ctrl_inst.latch_mem_inst.RAM\[55\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[44\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND net204 dig_ctrl_inst.latch_mem_inst.gclk\[44\] dig_ctrl_inst.latch_mem_inst.RAM\[44\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
X_2030_ VGND VDPWR VDPWR VGND _0686_ _0689_ _0688_ dig_ctrl_inst.latch_mem_inst.RAM\[39\]\[6\]
+ _0142_ _0687_ sky130_fd_sc_hd__a2111o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[33\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND net226 dig_ctrl_inst.latch_mem_inst.gclk\[33\] dig_ctrl_inst.latch_mem_inst.RAM\[33\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
X_1814_ VDPWR VGND VDPWR VGND net112 _0476_ dig_ctrl_inst.latch_mem_inst.RAM\[50\]\[3\]
+ net39 sky130_fd_sc_hd__and3_2
X_1745_ VDPWR VGND VDPWR VGND net112 _0408_ dig_ctrl_inst.latch_mem_inst.RAM\[18\]\[2\]
+ net60 sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[22\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND net242 dig_ctrl_inst.latch_mem_inst.gclk\[22\] dig_ctrl_inst.latch_mem_inst.RAM\[22\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
X_1676_ VGND VDPWR VDPWR VGND _0270_ _0340_ net261 _0027_ sky130_fd_sc_hd__mux2_1
X_2159_ VGND VDPWR VDPWR VGND _1039_ _0805_ net247 _0804_ sky130_fd_sc_hd__nand3_2
X_2228_ VDPWR VGND VDPWR VGND _0841_ _0262_ _0247_ _0872_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_39_Left_117 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.genblk1\[12\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[12\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[12\]._gclk clknet_leaf_19_clk sky130_fd_sc_hd__dlclkp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[59\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND net185 dig_ctrl_inst.latch_mem_inst.gclk\[59\] dig_ctrl_inst.latch_mem_inst.RAM\[59\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[10\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND net178 dig_ctrl_inst.latch_mem_inst.gclk\[10\] dig_ctrl_inst.latch_mem_inst.RAM\[10\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_48_Left_126 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_57_Left_135 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[48\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND net195 dig_ctrl_inst.latch_mem_inst.gclk\[48\] dig_ctrl_inst.latch_mem_inst.RAM\[48\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[4\].gen_latches\[0\].p_latch VGND VDPWR VDPWR
+ VGND net238 dig_ctrl_inst.latch_mem_inst.gclk\[4\] dig_ctrl_inst.latch_mem_inst.RAM\[4\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
X_1392_ VDPWR VGND VDPWR VGND net82 dig_ctrl_inst.latch_mem_inst.data_we\[26\] net146
+ net66 sky130_fd_sc_hd__and3_2
X_1530_ VGND VDPWR VDPWR VGND _0191_ _1104_ dig_ctrl_inst.cpu_inst.data\[1\] _0201_
+ sky130_fd_sc_hd__mux2_1
X_1461_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[62\] _0162_ net141
+ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_66_Left_144 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[37\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND net212 dig_ctrl_inst.latch_mem_inst.gclk\[37\] dig_ctrl_inst.latch_mem_inst.RAM\[37\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
X_2013_ VGND VDPWR VDPWR VGND _0672_ net116 dig_ctrl_inst.latch_mem_inst.RAM\[49\]\[6\]
+ net138 net37 sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_75_Left_153 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_15_clk VGND VDPWR VDPWR VGND clknet_leaf_15_clk clknet_1_0__leaf_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_60_338 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1728_ VGND VDPWR VDPWR VGND _0389_ _0392_ _0391_ dig_ctrl_inst.latch_mem_inst.RAM\[33\]\[1\]
+ _0136_ _0390_ sky130_fd_sc_hd__a2111o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[26\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND net231 dig_ctrl_inst.latch_mem_inst.gclk\[26\] dig_ctrl_inst.latch_mem_inst.RAM\[26\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_13_254 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_1659_ VGND VDPWR VDPWR VGND _0324_ net77 dig_ctrl_inst.latch_mem_inst.RAM\[61\]\[0\]
+ net121 net46 sky130_fd_sc_hd__and4_1
XFILLER_0_0_181 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_176 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_63_132 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
Xdig_ctrl_inst.latch_mem_inst.gen_words\[8\].gen_latches\[1\].p_latch VGND VDPWR VDPWR
+ VGND net231 dig_ctrl_inst.latch_mem_inst.gclk\[8\] dig_ctrl_inst.latch_mem_inst.RAM\[8\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
X_2562_ VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_data_o\[6\] net175 _0086_ clknet_leaf_3_clk
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_338 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_40_23 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2493_ VDPWR VGND VDPWR VGND dig_ctrl_inst.cpu_inst.port_o\[7\] clknet_leaf_6_clk
+ _0019_ sky130_fd_sc_hd__dfxtp_1
X_1513_ VGND VDPWR VDPWR VGND _0190_ dig_ctrl_inst.cpu_inst.port_o\[2\] net359 _0014_
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_4_clk VGND VDPWR VDPWR VGND clknet_leaf_4_clk clknet_1_1__leaf_clk sky130_fd_sc_hd__clkbuf_8
X_1375_ VDPWR VGND VDPWR VGND net121 _0122_ net137 net68 sky130_fd_sc_hd__and3_2
X_1444_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[53\] _0154_ net148
+ sky130_fd_sc_hd__and2_1
XFILLER_0_65_53 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[19\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND net240 dig_ctrl_inst.latch_mem_inst.gclk\[19\] dig_ctrl_inst.latch_mem_inst.RAM\[19\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_5_262 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
Xfanout72 VGND VDPWR VDPWR VGND _0115_ net72 sky130_fd_sc_hd__clkbuf_2
Xfanout94 VGND VDPWR VDPWR VGND net94 net96 sky130_fd_sc_hd__clkbuf_4
Xfanout83 VGND VDPWR VDPWR VGND net83 _1189_ sky130_fd_sc_hd__clkbuf_4
Xfanout61 VGND VDPWR VDPWR VGND net70 net61 sky130_fd_sc_hd__clkbuf_2
Xfanout50 VGND VDPWR VDPWR VGND net51 net50 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_19_35 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_19_57 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_1993_ VGND VDPWR VDPWR VGND _0652_ net77 dig_ctrl_inst.latch_mem_inst.RAM\[45\]\[6\]
+ net119 net57 sky130_fd_sc_hd__and4_1
XFILLER_0_27_132 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2545_ VGND VDPWR VDPWR VGND dig_ctrl_inst.mode_sync net168 net292 clknet_leaf_4_clk
+ sky130_fd_sc_hd__dfrtp_1
X_2614_ VDPWR VGND VDPWR VGND uio_out[6] net277 sky130_fd_sc_hd__buf_2
X_2476_ VGND VDPWR VDPWR VGND dig_ctrl_inst.synchronizer_port_ms_i_inst.pipe\[0\]
+ net175 net1 clknet_leaf_8_clk sky130_fd_sc_hd__dfrtp_1
X_1358_ VDPWR VGND VDPWR VGND net124 _1190_ net83 sky130_fd_sc_hd__and2_2
X_1427_ VDPWR VGND VDPWR VGND net71 dig_ctrl_inst.latch_mem_inst.data_we\[44\] net141
+ net48 sky130_fd_sc_hd__and3_2
X_1289_ VGND VDPWR VDPWR VGND _1056_ _1071_ _1131_ _1130_ sky130_fd_sc_hd__or3_2
XFILLER_0_33_113 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
Xclkload3 VGND VDPWR VDPWR VGND clkload3/Y clknet_leaf_12_clk sky130_fd_sc_hd__inv_16
Xfanout240 VDPWR VGND VDPWR VGND net240 net241 sky130_fd_sc_hd__buf_2
Xfanout251 VDPWR VGND VDPWR VGND net251 net252 sky130_fd_sc_hd__buf_2
Xfanout262 VDPWR VGND VDPWR VGND net262 net263 sky130_fd_sc_hd__buf_2
XFILLER_0_21_69 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2330_ VGND VDPWR VDPWR VGND _0970_ _0969_ _0968_ sky130_fd_sc_hd__nand2_1
X_2261_ VDPWR VGND VDPWR VGND dig_ctrl_inst.spi_data_o\[3\] _0183_ _0904_ dig_ctrl_inst.synchronizer_port_i_inst\[3\].out
+ _0824_ sky130_fd_sc_hd__a22o_1
X_2192_ VGND VDPWR VDPWR VGND net150 _0799_ _0790_ _0837_ sky130_fd_sc_hd__mux2_1
X_1212_ VDPWR VGND VDPWR VGND dig_ctrl_inst.cpu_inst.cpu_state\[1\] net245 dig_ctrl_inst.cpu_inst.cpu_state\[0\]
+ _1054_ sky130_fd_sc_hd__or3b_2
X_1976_ VDPWR VGND VDPWR VGND _0634_ _0632_ _0636_ _0633_ _0635_ sky130_fd_sc_hd__or4_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[63\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND net221 dig_ctrl_inst.latch_mem_inst.gclk\[63\] dig_ctrl_inst.latch_mem_inst.RAM\[63\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
X_2528_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[1\]\[0\] net156 _0054_
+ clknet_leaf_8_clk sky130_fd_sc_hd__dfrtp_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[17\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[17\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[17\]._gclk clknet_leaf_1_clk sky130_fd_sc_hd__dlclkp_1
XFILLER_0_30_149 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xhold15 VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_receiver_inst.synchronizer_spi_sclk.pipe\[0\]
+ net297 sky130_fd_sc_hd__dlygate4sd3_1
X_2459_ VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_receiver_inst.spi_cnt\[2\] net174
+ _0003_ clknet_leaf_5_clk sky130_fd_sc_hd__dfrtp_1
Xhold48 VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_miso_o net330 sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_data_i\[6\] net308 sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[0\]\[4\] net341 sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[3\]\[2\] net319 sky130_fd_sc_hd__dlygate4sd3_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[52\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND net239 dig_ctrl_inst.latch_mem_inst.gclk\[52\] dig_ctrl_inst.latch_mem_inst.RAM\[52\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_53_219 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[40\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND net179 dig_ctrl_inst.latch_mem_inst.gclk\[40\] dig_ctrl_inst.latch_mem_inst.RAM\[40\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
X_1830_ VDPWR VGND VDPWR VGND net133 _0492_ dig_ctrl_inst.latch_mem_inst.RAM\[16\]\[3\]
+ net59 sky130_fd_sc_hd__and3_2
X_1761_ VGND VDPWR VDPWR VGND _0421_ _0424_ _0423_ dig_ctrl_inst.latch_mem_inst.RAM\[46\]\[2\]
+ _0148_ _0422_ sky130_fd_sc_hd__a2111o_1
X_1692_ VGND VDPWR VDPWR VGND _0356_ net62 _1180_ dig_ctrl_inst.latch_mem_inst.RAM\[3\]\[1\]
+ dig_ctrl_inst.latch_mem_inst.RAM\[28\]\[1\] net72 sky130_fd_sc_hd__a32o_1
X_2313_ VGND VDPWR VDPWR VGND _0952_ _0953_ _0951_ sky130_fd_sc_hd__nor2_1
X_2244_ VGND VDPWR VDPWR VGND _0831_ _0887_ _0776_ sky130_fd_sc_hd__nor2_1
X_2175_ VDPWR VGND VDPWR VGND _0260_ _0814_ _0816_ _0821_ _0820_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_75_333 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_11_Left_89 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_7_165 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1959_ VGND VDPWR VDPWR VGND _0619_ net124 dig_ctrl_inst.latch_mem_inst.RAM\[1\]\[5\]
+ net138 net116 sky130_fd_sc_hd__and4_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[56\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND net229 dig_ctrl_inst.latch_mem_inst.gclk\[56\] dig_ctrl_inst.latch_mem_inst.RAM\[56\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
Xoutput16 VDPWR VGND VDPWR VGND port_ms_o[0] net16 sky130_fd_sc_hd__buf_2
Xoutput27 VDPWR VGND VDPWR VGND uo_out[2] net27 sky130_fd_sc_hd__buf_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[0\].gen_latches\[3\].p_latch VGND VDPWR VDPWR
+ VGND net213 dig_ctrl_inst.latch_mem_inst.gclk\[0\] dig_ctrl_inst.latch_mem_inst.RAM\[0\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
Xclkbuf_0_clk VGND VDPWR VDPWR VGND clknet_0_clk clk sky130_fd_sc_hd__clkbuf_16
Xdig_ctrl_inst.latch_mem_inst.gen_words\[33\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND net193 dig_ctrl_inst.latch_mem_inst.gclk\[33\] dig_ctrl_inst.latch_mem_inst.RAM\[33\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
X_1813_ VDPWR VGND VDPWR VGND net93 _0475_ dig_ctrl_inst.latch_mem_inst.RAM\[54\]\[3\]
+ net38 sky130_fd_sc_hd__and3_2
XFILLER_0_4_179 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_1744_ VDPWR VGND VDPWR VGND net93 _0407_ dig_ctrl_inst.latch_mem_inst.RAM\[54\]\[2\]
+ net40 sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[22\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND net210 dig_ctrl_inst.latch_mem_inst.gclk\[22\] dig_ctrl_inst.latch_mem_inst.RAM\[22\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_15_Right_15 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1675_ VDPWR VGND VDPWR VGND _0306_ _0340_ _0339_ _0279_ dig_ctrl_inst.latch_mem_inst.RAM\[0\]\[0\]
+ sky130_fd_sc_hd__o2bb2a_1
X_2089_ VDPWR VGND VDPWR VGND _0747_ _1184_ dig_ctrl_inst.latch_mem_inst.RAM\[1\]\[7\]
+ dig_ctrl_inst.latch_mem_inst.RAM\[7\]\[7\] _1175_ _0745_ sky130_fd_sc_hd__a221o_1
XFILLER_0_23_3 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_2227_ VGND VDPWR VDPWR VGND _0870_ _0815_ _0764_ _0871_ sky130_fd_sc_hd__mux2_1
X_2158_ VDPWR VGND VDPWR VGND _0804_ dig_ctrl_inst.cpu_inst.instr\[6\] dig_ctrl_inst.cpu_inst.instr\[7\]
+ sky130_fd_sc_hd__and2b_2
XPHY_EDGE_ROW_24_Right_24 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[11\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND net223 dig_ctrl_inst.latch_mem_inst.gclk\[11\] dig_ctrl_inst.latch_mem_inst.RAM\[11\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_33_Right_33 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[49\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND net243 dig_ctrl_inst.latch_mem_inst.gclk\[49\] dig_ctrl_inst.latch_mem_inst.RAM\[49\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_42_Right_42 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.genblk1\[42\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[42\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[42\]._gclk sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_51_Right_51 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[4\].gen_latches\[4\].p_latch VGND VDPWR VDPWR
+ VGND net210 dig_ctrl_inst.latch_mem_inst.gclk\[4\] dig_ctrl_inst.latch_mem_inst.RAM\[4\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
X_1391_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[25\] _0129_ net144
+ sky130_fd_sc_hd__and2_1
X_1460_ VDPWR VGND VDPWR VGND net75 _0162_ net114 net41 sky130_fd_sc_hd__and3_2
XPHY_EDGE_ROW_60_Right_60 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[37\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND net183 dig_ctrl_inst.latch_mem_inst.gclk\[37\] dig_ctrl_inst.latch_mem_inst.RAM\[37\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
X_2012_ VDPWR VGND VDPWR VGND net124 _0671_ dig_ctrl_inst.latch_mem_inst.RAM\[12\]\[6\]
+ net71 sky130_fd_sc_hd__and3_2
X_1727_ VDPWR VGND VDPWR VGND net135 _0391_ dig_ctrl_inst.latch_mem_inst.RAM\[16\]\[1\]
+ net65 sky130_fd_sc_hd__and3_2
X_1658_ VDPWR VGND VDPWR VGND net74 _0323_ dig_ctrl_inst.latch_mem_inst.RAM\[44\]\[0\]
+ net56 sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[26\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND net202 dig_ctrl_inst.latch_mem_inst.gclk\[26\] dig_ctrl_inst.latch_mem_inst.RAM\[26\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_0_193 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1589_ VGND VDPWR VDPWR VGND _0255_ _0172_ _0221_ sky130_fd_sc_hd__nand2b_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[15\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND net215 dig_ctrl_inst.latch_mem_inst.gclk\[15\] dig_ctrl_inst.latch_mem_inst.RAM\[15\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_48_141 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_14_Left_92 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_39_141 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
Xdig_ctrl_inst.latch_mem_inst.gen_words\[8\].gen_latches\[5\].p_latch VGND VDPWR VDPWR
+ VGND net195 dig_ctrl_inst.latch_mem_inst.gclk\[8\] dig_ctrl_inst.latch_mem_inst.RAM\[8\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
X_2492_ VDPWR VGND VDPWR VGND dig_ctrl_inst.cpu_inst.port_o\[6\] clknet_leaf_5_clk
+ _0018_ sky130_fd_sc_hd__dfxtp_1
X_1512_ VGND VDPWR VDPWR VGND _0190_ dig_ctrl_inst.cpu_inst.port_o\[1\] dig_ctrl_inst.cpu_inst.regs\[0\]\[1\]
+ _0013_ sky130_fd_sc_hd__mux2_1
X_2561_ VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_data_o\[5\] net175 _0085_ clknet_leaf_3_clk
+ sky130_fd_sc_hd__dfrtp_1
X_1443_ VDPWR VGND VDPWR VGND net102 _0154_ net119 net43 sky130_fd_sc_hd__and3_2
X_1374_ VDPWR VGND VDPWR VGND net141 dig_ctrl_inst.latch_mem_inst.data_we\[16\] net133
+ net61 sky130_fd_sc_hd__and3_2
XFILLER_0_4_24 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.genblk1\[1\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[1\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[1\]._gclk clknet_leaf_15_clk sky130_fd_sc_hd__dlclkp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[19\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND net205 dig_ctrl_inst.latch_mem_inst.gclk\[19\] dig_ctrl_inst.latch_mem_inst.RAM\[19\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
Xfanout73 VDPWR VGND VDPWR VGND net73 _0115_ sky130_fd_sc_hd__buf_2
Xfanout51 VGND VDPWR VDPWR VGND net52 net51 sky130_fd_sc_hd__clkbuf_2
Xdig_ctrl_inst.latch_mem_inst.genblk1\[24\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[24\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[24\]._gclk clknet_leaf_13_clk sky130_fd_sc_hd__dlclkp_1
Xfanout40 VGND VDPWR VDPWR VGND net40 net42 sky130_fd_sc_hd__buf_1
Xfanout62 VDPWR VGND VDPWR VGND net62 net70 sky130_fd_sc_hd__buf_2
Xfanout95 VGND VDPWR VDPWR VGND net96 net95 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_51_158 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_24_339 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xfanout84 VDPWR VGND VDPWR VGND net84 net87 sky130_fd_sc_hd__buf_2
X_2602__279 VGND VDPWR VDPWR VGND _2602__279/LO net279 sky130_fd_sc_hd__conb_1
X_1992_ VDPWR VGND VDPWR VGND net128 _0651_ dig_ctrl_inst.latch_mem_inst.RAM\[6\]\[6\]
+ net94 sky130_fd_sc_hd__and3_2
Xclkload10 VGND VDPWR VDPWR VGND clkload10/Y clknet_leaf_2_clk sky130_fd_sc_hd__clkinv_16
XFILLER_0_42_136 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2475_ VGND VDPWR VDPWR VGND dig_ctrl_inst.synchronizer_port_i_inst\[0\].out net170
+ net300 clknet_leaf_5_clk sky130_fd_sc_hd__dfrtp_1
X_2544_ VGND VDPWR VDPWR VGND dig_ctrl_inst.synchronizer_mode_i_inst.pipe\[0\] net168
+ net14 clknet_leaf_4_clk sky130_fd_sc_hd__dfrtp_1
X_2613_ VDPWR VGND VDPWR VGND uio_out[5] net276 sky130_fd_sc_hd__buf_2
X_1357_ VDPWR VGND VDPWR VGND _1189_ _1139_ _1122_ _1106_ _1090_ _1052_ sky130_fd_sc_hd__o2111a_1
X_1288_ VGND VDPWR VDPWR VGND _1063_ _1125_ _1126_ _1127_ _1130_ _1128_ sky130_fd_sc_hd__o41ai_2
X_1426_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[43\] _0146_ net143
+ sky130_fd_sc_hd__and2_1
XFILLER_0_33_169 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xclkload4 VGND VDPWR VDPWR VGND clkload4/Y clknet_leaf_13_clk sky130_fd_sc_hd__clkinv_1
XFILLER_0_18_166 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xfanout241 VGND VDPWR VDPWR VGND net244 net241 sky130_fd_sc_hd__clkbuf_2
Xdig_ctrl_inst.latch_mem_inst.genblk1\[35\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[35\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[35\]._gclk sky130_fd_sc_hd__clkbuf_4
Xfanout230 VGND VDPWR VDPWR VGND net290 net230 sky130_fd_sc_hd__clkbuf_2
Xfanout252 VDPWR VGND VDPWR VGND dig_ctrl_inst.cpu_inst.arg1\[1\] net252 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout263 VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.arg0\[0\] net263 sky130_fd_sc_hd__clkbuf_2
X_2191_ VGND VDPWR VDPWR VGND _0835_ _0836_ _0795_ sky130_fd_sc_hd__nor2_1
X_1211_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.cpu_state\[1\] dig_ctrl_inst.cpu_inst.cpu_state\[0\]
+ net245 _1053_ sky130_fd_sc_hd__nor3b_4
X_2260_ VGND VDPWR VDPWR VGND _0877_ _0903_ _1120_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_1_69 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1975_ VGND VDPWR VDPWR VGND _0594_ _0635_ _0604_ dig_ctrl_inst.latch_mem_inst.RAM\[33\]\[5\]
+ _0136_ _0601_ sky130_fd_sc_hd__a2111o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[63\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND net189 dig_ctrl_inst.latch_mem_inst.gclk\[63\] dig_ctrl_inst.latch_mem_inst.RAM\[63\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_11_70 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_15_169 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2458_ VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_receiver_inst.spi_cnt\[1\] net172
+ _0002_ clknet_leaf_5_clk sky130_fd_sc_hd__dfrtp_1
Xhold27 VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_data_i\[5\] net309 sky130_fd_sc_hd__dlygate4sd3_1
Xhold16 VGND VDPWR VDPWR VGND dig_ctrl_inst.synchronizer_port_i_inst\[3\].pipe\[0\]
+ net298 sky130_fd_sc_hd__dlygate4sd3_1
X_1409_ VGND VDPWR VDPWR VGND net137 net108 net57 _0138_ sky130_fd_sc_hd__and3_4
X_2527_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[0\]\[7\] net156 _0053_
+ clknet_leaf_8_clk sky130_fd_sc_hd__dfrtp_2
Xhold38 VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[2\]\[2\] net320 sky130_fd_sc_hd__dlygate4sd3_1
X_2389_ VGND VDPWR VDPWR VGND _1003_ _1001_ net334 _0077_ sky130_fd_sc_hd__mux2_1
Xhold49 VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[2\]\[4\] net331 sky130_fd_sc_hd__dlygate4sd3_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[52\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND net209 dig_ctrl_inst.latch_mem_inst.gclk\[52\] dig_ctrl_inst.latch_mem_inst.RAM\[52\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[41\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND net220 dig_ctrl_inst.latch_mem_inst.gclk\[41\] dig_ctrl_inst.latch_mem_inst.RAM\[41\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[30\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND net240 dig_ctrl_inst.latch_mem_inst.gclk\[30\] dig_ctrl_inst.latch_mem_inst.RAM\[30\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
X_1691_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[19\]\[1\] _0124_ _0355_
+ dig_ctrl_inst.latch_mem_inst.RAM\[53\]\[1\] _0154_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_317 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1760_ VDPWR VGND VDPWR VGND net83 _0423_ dig_ctrl_inst.latch_mem_inst.RAM\[58\]\[2\]
+ net38 sky130_fd_sc_hd__and3_2
XPHY_EDGE_ROW_2_Left_80 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2312_ VDPWR VGND VDPWR VGND _0952_ _0930_ _0231_ _0932_ sky130_fd_sc_hd__a21boi_1
X_2615__278 VGND VDPWR VDPWR VGND net278 _2615__278/HI sky130_fd_sc_hd__conb_1
X_2243_ VGND VDPWR VDPWR VGND _0797_ _0885_ _0886_ _0884_ sky130_fd_sc_hd__or3b_1
X_2174_ VGND VDPWR VDPWR VGND _0817_ _0820_ _0819_ sky130_fd_sc_hd__or2_1
Xoutput17 VDPWR VGND VDPWR VGND port_ms_o[1] net17 sky130_fd_sc_hd__buf_2
X_1958_ VGND VDPWR VDPWR VGND _0618_ net90 dig_ctrl_inst.latch_mem_inst.RAM\[59\]\[5\]
+ net108 net46 sky130_fd_sc_hd__and4_1
Xoutput28 VDPWR VGND VDPWR VGND uo_out[3] net28 sky130_fd_sc_hd__buf_2
X_1889_ VDPWR VGND VDPWR VGND _0550_ _0149_ dig_ctrl_inst.latch_mem_inst.RAM\[27\]\[4\]
+ dig_ctrl_inst.latch_mem_inst.RAM\[47\]\[4\] _0130_ _0549_ sky130_fd_sc_hd__a221o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[56\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND net199 dig_ctrl_inst.latch_mem_inst.gclk\[56\] dig_ctrl_inst.latch_mem_inst.RAM\[56\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[45\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND net218 dig_ctrl_inst.latch_mem_inst.gclk\[45\] dig_ctrl_inst.latch_mem_inst.RAM\[45\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_34_231 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[34\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND net230 dig_ctrl_inst.latch_mem_inst.gclk\[34\] dig_ctrl_inst.latch_mem_inst.RAM\[34\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[0\].gen_latches\[7\].p_latch VGND VDPWR VDPWR
+ VGND net180 dig_ctrl_inst.latch_mem_inst.gclk\[0\] dig_ctrl_inst.latch_mem_inst.RAM\[0\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
X_1743_ VDPWR VGND VDPWR VGND _0403_ _0406_ _0404_ _0405_ sky130_fd_sc_hd__or3_1
X_1812_ VDPWR VGND VDPWR VGND net71 _0474_ dig_ctrl_inst.latch_mem_inst.RAM\[60\]\[3\]
+ net38 sky130_fd_sc_hd__and3_2
X_1674_ VGND VDPWR VDPWR VGND _0338_ _0321_ _0277_ _0271_ _0339_ sky130_fd_sc_hd__o211a_1
XFILLER_0_68_76 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2226_ VDPWR VGND VDPWR VGND _0870_ _0869_ _0868_ sky130_fd_sc_hd__and2_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[6\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[6\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[6\]._gclk clknet_leaf_13_clk sky130_fd_sc_hd__dlclkp_1
X_2088_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[30\]\[7\] _0132_ _0746_
+ dig_ctrl_inst.latch_mem_inst.RAM\[63\]\[7\] _0163_ sky130_fd_sc_hd__a22o_1
X_2157_ VGND VDPWR VDPWR VGND _0803_ _0787_ _0802_ _1129_ _1113_ sky130_fd_sc_hd__a211o_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[29\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[29\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[29\]._gclk clknet_leaf_15_clk sky130_fd_sc_hd__dlclkp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[11\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND net190 dig_ctrl_inst.latch_mem_inst.gclk\[11\] dig_ctrl_inst.latch_mem_inst.RAM\[11\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[28\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[28\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[28\]._gclk sky130_fd_sc_hd__clkbuf_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[49\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND net209 dig_ctrl_inst.latch_mem_inst.gclk\[49\] dig_ctrl_inst.latch_mem_inst.RAM\[49\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[38\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND net225 dig_ctrl_inst.latch_mem_inst.gclk\[38\] dig_ctrl_inst.latch_mem_inst.RAM\[38\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_1_139 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.genblk1\[31\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[31\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[31\]._gclk clknet_leaf_17_clk sky130_fd_sc_hd__dlclkp_1
X_1390_ VDPWR VGND VDPWR VGND net89 _0129_ net117 net60 sky130_fd_sc_hd__and3_2
XFILLER_0_49_109 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[27\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND net236 dig_ctrl_inst.latch_mem_inst.gclk\[27\] dig_ctrl_inst.latch_mem_inst.RAM\[27\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
X_2011_ VDPWR VGND VDPWR VGND net93 _0670_ dig_ctrl_inst.latch_mem_inst.RAM\[54\]\[6\]
+ net37 sky130_fd_sc_hd__and3_2
X_1726_ VDPWR VGND VDPWR VGND net127 _0390_ dig_ctrl_inst.latch_mem_inst.RAM\[4\]\[1\]
+ net100 sky130_fd_sc_hd__and3_2
X_1657_ VGND VDPWR VDPWR VGND _0322_ net107 dig_ctrl_inst.latch_mem_inst.RAM\[7\]\[0\]
+ net129 net101 sky130_fd_sc_hd__and4_1
X_1588_ VGND VDPWR VDPWR VGND _0168_ _0227_ _0254_ _0224_ sky130_fd_sc_hd__or3b_1
X_2209_ VDPWR VGND VDPWR VGND dig_ctrl_inst.spi_data_o\[1\] _0183_ _0854_ dig_ctrl_inst.synchronizer_port_i_inst\[1\].out
+ _0824_ sky130_fd_sc_hd__a22o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[15\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND net179 dig_ctrl_inst.latch_mem_inst.gclk\[15\] dig_ctrl_inst.latch_mem_inst.RAM\[15\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[9\].gen_latches\[0\].p_latch VGND VDPWR VDPWR
+ VGND net238 dig_ctrl_inst.latch_mem_inst.gclk\[9\] dig_ctrl_inst.latch_mem_inst.RAM\[9\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_5_3 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_39_153 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_27_337 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2560_ VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_data_o\[4\] net175 _0084_ clknet_leaf_9_clk
+ sky130_fd_sc_hd__dfrtp_1
X_1511_ VGND VDPWR VDPWR VGND _0190_ dig_ctrl_inst.cpu_inst.port_o\[0\] dig_ctrl_inst.cpu_inst.regs\[0\]\[0\]
+ _0012_ sky130_fd_sc_hd__mux2_1
X_2491_ VDPWR VGND VDPWR VGND dig_ctrl_inst.cpu_inst.port_o\[5\] clknet_leaf_6_clk
+ _0017_ sky130_fd_sc_hd__dfxtp_1
X_1442_ VDPWR VGND VDPWR VGND net98 dig_ctrl_inst.latch_mem_inst.data_we\[52\] net147
+ net46 sky130_fd_sc_hd__and3_2
X_1373_ VDPWR VGND VDPWR VGND _0121_ net65 net135 sky130_fd_sc_hd__and2_1
X_1709_ VGND VDPWR VDPWR VGND _0370_ _0373_ _0372_ dig_ctrl_inst.latch_mem_inst.RAM\[15\]\[1\]
+ _0119_ _0371_ sky130_fd_sc_hd__a2111o_1
Xfanout96 VDPWR VGND VDPWR VGND net96 _1183_ sky130_fd_sc_hd__buf_2
Xfanout74 VGND VDPWR VDPWR VGND net74 _0115_ sky130_fd_sc_hd__buf_1
Xfanout63 VGND VDPWR VDPWR VGND net64 net63 sky130_fd_sc_hd__clkbuf_2
Xfanout41 VDPWR VGND VDPWR VGND net41 net42 sky130_fd_sc_hd__buf_2
Xfanout52 VDPWR VGND VDPWR VGND net52 _0134_ sky130_fd_sc_hd__buf_2
Xfanout85 VGND VDPWR VDPWR VGND net87 net85 sky130_fd_sc_hd__clkbuf_2
Xdig_ctrl_inst.latch_mem_inst.genblk1\[8\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[8\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[8\]._gclk sky130_fd_sc_hd__clkbuf_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[60\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND net236 dig_ctrl_inst.latch_mem_inst.gclk\[60\] dig_ctrl_inst.latch_mem_inst.RAM\[60\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
Xclkload11 VGND VDPWR VDPWR VGND clknet_leaf_3_clk clkload11/Y sky130_fd_sc_hd__inv_12
X_2612_ VDPWR VGND VDPWR VGND uio_out[4] net275 sky130_fd_sc_hd__buf_2
XFILLER_0_42_104 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
X_1991_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[1\]\[6\] _1175_ _0650_
+ dig_ctrl_inst.latch_mem_inst.RAM\[62\]\[6\] _0162_ sky130_fd_sc_hd__a22o_1
X_2474_ VGND VDPWR VDPWR VGND dig_ctrl_inst.synchronizer_port_i_inst\[0\].pipe\[0\]
+ net169 net3 clknet_leaf_4_clk sky130_fd_sc_hd__dfrtp_1
X_2543_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[2\]\[7\] net153 _0069_
+ clknet_leaf_11_clk sky130_fd_sc_hd__dfrtp_1
X_1425_ VDPWR VGND VDPWR VGND net89 _0146_ net104 net50 sky130_fd_sc_hd__and3_2
X_1287_ VGND VDPWR VDPWR VGND _1063_ _1125_ _1126_ _1127_ _1128_ _1129_ sky130_fd_sc_hd__o41a_4
X_1356_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[9\] _1188_ net141
+ sky130_fd_sc_hd__and2_1
Xclkload5 VGND VDPWR VDPWR VGND clkload5/Y clknet_leaf_14_clk sky130_fd_sc_hd__inv_16
Xfanout264 VGND VDPWR VDPWR VGND net264 net265 sky130_fd_sc_hd__clkbuf_4
Xfanout242 VDPWR VGND VDPWR VGND net242 net243 sky130_fd_sc_hd__buf_2
Xfanout231 VGND VDPWR VDPWR VGND net232 net231 sky130_fd_sc_hd__clkbuf_2
Xfanout220 VGND VDPWR VDPWR VGND net221 net220 sky130_fd_sc_hd__clkbuf_2
Xfanout253 VDPWR VGND VDPWR VGND net253 net254 sky130_fd_sc_hd__buf_2
XFILLER_0_49_281 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_1210_ VGND VDPWR VDPWR VGND _1041_ _1052_ dig_ctrl_inst.spi_addr\[0\] sky130_fd_sc_hd__nor2_2
X_2190_ VGND VDPWR VDPWR VGND net149 _0790_ _0788_ _0835_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_15 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_1974_ VGND VDPWR VDPWR VGND _0580_ _0634_ _0612_ dig_ctrl_inst.latch_mem_inst.RAM\[61\]\[5\]
+ _0161_ _0603_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_7_337 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2457_ VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_receiver_inst.spi_cnt\[0\] net172
+ _0001_ clknet_leaf_5_clk sky130_fd_sc_hd__dfrtp_4
X_2388_ VGND VDPWR VDPWR VGND _1003_ _0999_ net345 _0076_ sky130_fd_sc_hd__mux2_1
Xhold17 VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_receiver_inst.synchronizer_spi_mosi.pipe\[0\]
+ net299 sky130_fd_sc_hd__dlygate4sd3_1
Xhold39 VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[2\]\[5\] net321 sky130_fd_sc_hd__dlygate4sd3_1
X_2526_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[0\]\[6\] net157 _0052_
+ clknet_leaf_9_clk sky130_fd_sc_hd__dfrtp_1
Xhold28 VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.prev_state\[2\] net310 sky130_fd_sc_hd__dlygate4sd3_1
X_1408_ VDPWR VGND VDPWR VGND net111 dig_ctrl_inst.latch_mem_inst.data_we\[34\] net141
+ net48 sky130_fd_sc_hd__and3_2
X_1339_ VDPWR VGND VDPWR VGND net143 dig_ctrl_inst.latch_mem_inst.data_we\[2\] net125
+ net112 sky130_fd_sc_hd__and3_2
XFILLER_0_21_118 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
Xdig_ctrl_inst.latch_mem_inst.gen_words\[41\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND net188 dig_ctrl_inst.latch_mem_inst.gclk\[41\] dig_ctrl_inst.latch_mem_inst.RAM\[41\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[36\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[36\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[36\]._gclk clknet_leaf_4_clk sky130_fd_sc_hd__dlclkp_1
XFILLER_0_16_38 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[30\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND net209 dig_ctrl_inst.latch_mem_inst.gclk\[30\] dig_ctrl_inst.latch_mem_inst.RAM\[30\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
X_1690_ VGND VDPWR VDPWR VGND _0351_ _0354_ _0353_ dig_ctrl_inst.latch_mem_inst.RAM\[21\]\[1\]
+ _0126_ _0352_ sky130_fd_sc_hd__a2111o_1
X_2242_ VGND VDPWR VDPWR VGND _0830_ _0885_ _0834_ _0782_ _0776_ sky130_fd_sc_hd__o22a_1
X_2311_ VGND VDPWR VDPWR VGND _0231_ _0930_ _0951_ _0932_ sky130_fd_sc_hd__and3b_1
X_2173_ VGND VDPWR VDPWR VGND _1039_ _0819_ _0774_ net247 sky130_fd_sc_hd__and3b_2
X_1957_ VGND VDPWR VDPWR VGND _0617_ net76 dig_ctrl_inst.latch_mem_inst.RAM\[31\]\[5\]
+ net106 net64 sky130_fd_sc_hd__and4_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[57\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND net242 dig_ctrl_inst.latch_mem_inst.gclk\[57\] dig_ctrl_inst.latch_mem_inst.RAM\[57\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_22_81 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xoutput18 VDPWR VGND VDPWR VGND port_ms_o[2] net18 sky130_fd_sc_hd__buf_2
Xoutput29 VDPWR VGND VDPWR VGND uo_out[4] net29 sky130_fd_sc_hd__buf_2
X_1888_ VGND VDPWR VDPWR VGND _0549_ net64 dig_ctrl_inst.latch_mem_inst.RAM\[16\]\[4\]
+ _0121_ dig_ctrl_inst.latch_mem_inst.RAM\[26\]\[4\] net81 sky130_fd_sc_hd__a32o_1
X_2509_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.data\[0\] net153 _0035_ clknet_leaf_10_clk
+ sky130_fd_sc_hd__dfrtp_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[45\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND net182 dig_ctrl_inst.latch_mem_inst.gclk\[45\] dig_ctrl_inst.latch_mem_inst.RAM\[45\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[1\].gen_latches\[2\].p_latch VGND VDPWR VDPWR
+ VGND net220 dig_ctrl_inst.latch_mem_inst.gclk\[1\] dig_ctrl_inst.latch_mem_inst.RAM\[1\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[34\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND net195 dig_ctrl_inst.latch_mem_inst.gclk\[34\] dig_ctrl_inst.latch_mem_inst.RAM\[34\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
X_1811_ VGND VDPWR VDPWR VGND _0473_ net92 dig_ctrl_inst.latch_mem_inst.RAM\[41\]\[3\]
+ net118 net53 sky130_fd_sc_hd__and4_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[23\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND net217 dig_ctrl_inst.latch_mem_inst.gclk\[23\] dig_ctrl_inst.latch_mem_inst.RAM\[23\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
X_1742_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[42\]\[2\] _0145_ _0405_
+ dig_ctrl_inst.latch_mem_inst.RAM\[59\]\[2\] _0159_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_321 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_1673_ VGND VDPWR VDPWR VGND _0337_ _0333_ _0338_ _0325_ _0329_ sky130_fd_sc_hd__nor4_1
XFILLER_0_7_69 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2225_ VGND VDPWR VDPWR VGND _0869_ _0850_ net160 sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_18_clk VGND VDPWR VDPWR VGND clknet_leaf_18_clk clknet_1_1__leaf_clk
+ sky130_fd_sc_hd__clkbuf_8
Xdig_ctrl_inst.latch_mem_inst.gen_words\[12\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND net232 dig_ctrl_inst.latch_mem_inst.gclk\[12\] dig_ctrl_inst.latch_mem_inst.RAM\[12\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
X_2087_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[16\]\[7\] _0121_ _0745_
+ dig_ctrl_inst.latch_mem_inst.RAM\[61\]\[7\] _0161_ sky130_fd_sc_hd__a22o_1
X_2156_ VGND VDPWR VDPWR VGND _0802_ _0776_ _0801_ _0792_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_5_Right_5 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[5\].gen_latches\[3\].p_latch VGND VDPWR VDPWR
+ VGND net215 dig_ctrl_inst.latch_mem_inst.gclk\[5\] dig_ctrl_inst.latch_mem_inst.RAM\[5\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_26_Left_104 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[38\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND net189 dig_ctrl_inst.latch_mem_inst.gclk\[38\] dig_ctrl_inst.latch_mem_inst.RAM\[38\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
X_2010_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[2\]\[6\] _1178_ _0669_
+ dig_ctrl_inst.latch_mem_inst.RAM\[32\]\[6\] _0135_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_35_Left_113 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1725_ VGND VDPWR VDPWR VGND _0389_ net91 dig_ctrl_inst.latch_mem_inst.RAM\[25\]\[1\]
+ net118 net65 sky130_fd_sc_hd__and4_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[27\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND net209 dig_ctrl_inst.latch_mem_inst.gclk\[27\] dig_ctrl_inst.latch_mem_inst.RAM\[27\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_44_Left_122 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_7_clk VGND VDPWR VDPWR VGND clknet_leaf_7_clk clknet_1_1__leaf_clk sky130_fd_sc_hd__clkbuf_8
X_1656_ VGND VDPWR VDPWR VGND _0320_ _0316_ _0321_ _0310_ _0314_ sky130_fd_sc_hd__nor4_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[16\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND net220 dig_ctrl_inst.latch_mem_inst.gclk\[16\] dig_ctrl_inst.latch_mem_inst.RAM\[16\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
X_1587_ VGND VDPWR VDPWR VGND _0251_ _0232_ _0250_ _0252_ _0253_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_53_Left_131 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2139_ VDPWR VGND VDPWR VGND _0785_ _0777_ _0221_ sky130_fd_sc_hd__and2_1
X_2208_ VDPWR VGND VDPWR VGND _0843_ _0853_ _0848_ _0852_ sky130_fd_sc_hd__or3_1
XFILLER_0_48_154 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_62_Left_140 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_8_284 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_24_49 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[9\].gen_latches\[4\].p_latch VGND VDPWR VDPWR
+ VGND net204 dig_ctrl_inst.latch_mem_inst.gclk\[9\] dig_ctrl_inst.latch_mem_inst.RAM\[9\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_54_157 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2490_ VDPWR VGND VDPWR VGND dig_ctrl_inst.cpu_inst.port_o\[4\] clknet_leaf_6_clk
+ _0016_ sky130_fd_sc_hd__dfxtp_1
X_1510_ VDPWR VGND VDPWR VGND _1051_ _1067_ dig_ctrl_inst.cpu_inst.skip _0186_ _0190_
+ sky130_fd_sc_hd__or4_4
X_1441_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[51\] _0153_ net148
+ sky130_fd_sc_hd__and2_1
X_1372_ VGND VDPWR VDPWR VGND _0120_ _1156_ _1170_ sky130_fd_sc_hd__and2b_1
XFILLER_0_18_305 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_60_149 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_76_3 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1708_ VGND VDPWR VDPWR VGND _0372_ net77 dig_ctrl_inst.latch_mem_inst.RAM\[30\]\[1\]
+ net114 net65 sky130_fd_sc_hd__and4_1
X_1639_ VGND VDPWR VDPWR VGND _0301_ _0304_ _0303_ dig_ctrl_inst.latch_mem_inst.RAM\[29\]\[0\]
+ _0131_ _0302_ sky130_fd_sc_hd__a2111o_1
Xfanout53 VDPWR VGND VDPWR VGND net53 net54 sky130_fd_sc_hd__buf_2
Xfanout86 VDPWR VGND VDPWR VGND net86 net87 sky130_fd_sc_hd__buf_2
Xfanout64 VDPWR VGND VDPWR VGND net65 net64 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout75 VDPWR VGND VDPWR VGND net75 net76 sky130_fd_sc_hd__buf_2
XFILLER_0_36_124 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
Xfanout42 VGND VDPWR VDPWR VGND _0150_ net42 sky130_fd_sc_hd__clkbuf_2
Xfanout97 VDPWR VGND VDPWR VGND net97 _1182_ sky130_fd_sc_hd__buf_2
XFILLER_0_27_102 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_1990_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[40\]\[6\] _0143_ _0649_
+ dig_ctrl_inst.latch_mem_inst.RAM\[43\]\[6\] _0146_ sky130_fd_sc_hd__a22o_1
Xclkload12 VDPWR VGND VDPWR VGND clknet_leaf_5_clk clkload12/Y sky130_fd_sc_hd__clkinvlp_4
X_2542_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[2\]\[6\] net157 _0068_
+ clknet_leaf_7_clk sky130_fd_sc_hd__dfrtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[60\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND net207 dig_ctrl_inst.latch_mem_inst.gclk\[60\] dig_ctrl_inst.latch_mem_inst.RAM\[60\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
X_2611_ VDPWR VGND VDPWR VGND uio_out[3] net274 sky130_fd_sc_hd__buf_2
Xdig_ctrl_inst.latch_mem_inst.genblk1\[43\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[43\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[43\]._gclk clknet_leaf_15_clk sky130_fd_sc_hd__dlclkp_1
X_2473_ VGND VDPWR VDPWR VGND dig_ctrl_inst.synchronizer_port_i_inst\[1\].out net169
+ net302 clknet_leaf_5_clk sky130_fd_sc_hd__dfrtp_1
X_1424_ VDPWR VGND VDPWR VGND net82 dig_ctrl_inst.latch_mem_inst.data_we\[42\] net145
+ net55 sky130_fd_sc_hd__and3_2
X_1355_ VDPWR VGND VDPWR VGND net116 _1188_ net124 net88 sky130_fd_sc_hd__and3_2
X_1286_ VDPWR VGND VDPWR VGND net254 _1128_ net250 dig_ctrl_inst.cpu_inst.regs\[0\]\[2\]
+ sky130_fd_sc_hd__or3_1
Xclkload6 VGND VDPWR VDPWR VGND clknet_leaf_15_clk clkload6/Y sky130_fd_sc_hd__inv_12
Xfanout265 VDPWR VGND VDPWR VGND net265 net266 sky130_fd_sc_hd__buf_2
Xfanout232 VGND VDPWR VDPWR VGND net290 net232 sky130_fd_sc_hd__clkbuf_2
Xfanout243 VDPWR VGND VDPWR VGND net243 net244 sky130_fd_sc_hd__buf_2
Xfanout210 VGND VDPWR VDPWR VGND net283 net210 sky130_fd_sc_hd__clkbuf_2
Xfanout221 VGND VDPWR VDPWR VGND net221 net222 sky130_fd_sc_hd__buf_1
Xfanout254 VGND VDPWR VDPWR VGND net256 net254 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_5_80 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_46_25 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1973_ VGND VDPWR VDPWR VGND _0584_ _0633_ _0618_ dig_ctrl_inst.latch_mem_inst.RAM\[23\]\[5\]
+ _0128_ _0614_ sky130_fd_sc_hd__a2111o_1
X_2525_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[0\]\[5\] net157 _0051_
+ clknet_leaf_7_clk sky130_fd_sc_hd__dfrtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[53\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND net212 dig_ctrl_inst.latch_mem_inst.gclk\[53\] dig_ctrl_inst.latch_mem_inst.RAM\[53\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_39_3 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2456_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.rst_ni net282 net2 sky130_fd_sc_hd__dfxtp_1
Xhold29 VGND VDPWR VDPWR VGND net23 net311 sky130_fd_sc_hd__dlygate4sd3_1
X_2387_ VGND VDPWR VDPWR VGND _1003_ _0998_ net312 _0075_ sky130_fd_sc_hd__mux2_1
Xhold18 VGND VDPWR VDPWR VGND dig_ctrl_inst.synchronizer_port_i_inst\[0\].pipe\[0\]
+ net300 sky130_fd_sc_hd__dlygate4sd3_1
X_1338_ VDPWR VGND VDPWR VGND net124 _1178_ net111 sky130_fd_sc_hd__and2_2
X_1407_ VDPWR VGND VDPWR VGND _0137_ net48 net111 sky130_fd_sc_hd__and2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[42\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND net231 dig_ctrl_inst.latch_mem_inst.gclk\[42\] dig_ctrl_inst.latch_mem_inst.RAM\[42\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_36_91 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_1269_ VGND VDPWR VDPWR VGND _1111_ net254 dig_ctrl_inst.cpu_inst.regs\[2\]\[3\]
+ sky130_fd_sc_hd__nand2b_1
XFILLER_0_21_108 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_69_333 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.genblk1\[31\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[31\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[31\]._gclk sky130_fd_sc_hd__clkbuf_4
X_2310_ VDPWR VGND VDPWR VGND _0051_ _0950_ _0771_ _0946_ _0772_ net343 sky130_fd_sc_hd__o32a_1
XFILLER_0_57_57 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2172_ VGND VDPWR VDPWR VGND _0818_ _0773_ _0804_ sky130_fd_sc_hd__nand2b_1
X_2241_ VGND VDPWR VDPWR VGND _0857_ _0883_ _0884_ _0835_ _0795_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_43_233 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
X_1887_ VDPWR VGND VDPWR VGND _0546_ _0544_ _0548_ _0545_ _0547_ sky130_fd_sc_hd__or4_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[57\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND net208 dig_ctrl_inst.latch_mem_inst.gclk\[57\] dig_ctrl_inst.latch_mem_inst.RAM\[57\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
X_1956_ VGND VDPWR VDPWR VGND _0616_ net88 dig_ctrl_inst.latch_mem_inst.RAM\[41\]\[5\]
+ net116 net48 sky130_fd_sc_hd__and4_1
Xoutput19 VDPWR VGND VDPWR VGND port_ms_o[3] net19 sky130_fd_sc_hd__buf_2
X_2508_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.instr\[7\] net151 _0034_ clknet_leaf_13_clk
+ sky130_fd_sc_hd__dfrtp_4
X_2439_ VGND VDPWR VDPWR VGND _1024_ _1023_ dig_ctrl_inst.spi_addr\[0\] sky130_fd_sc_hd__nand2_1
XFILLER_0_47_90 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[46\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND net219 dig_ctrl_inst.latch_mem_inst.gclk\[46\] dig_ctrl_inst.latch_mem_inst.RAM\[46\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[35\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND net238 dig_ctrl_inst.latch_mem_inst.gclk\[35\] dig_ctrl_inst.latch_mem_inst.RAM\[35\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[1\].gen_latches\[6\].p_latch VGND VDPWR VDPWR
+ VGND net187 dig_ctrl_inst.latch_mem_inst.gclk\[1\] dig_ctrl_inst.latch_mem_inst.RAM\[1\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
X_1810_ VDPWR VGND VDPWR VGND net83 _0472_ dig_ctrl_inst.latch_mem_inst.RAM\[42\]\[3\]
+ net50 sky130_fd_sc_hd__and3_2
X_1741_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[3\]\[2\] _1180_ _0404_
+ dig_ctrl_inst.latch_mem_inst.RAM\[10\]\[2\] _1190_ sky130_fd_sc_hd__a22o_1
X_1672_ VGND VDPWR VDPWR VGND _0334_ _0337_ _0336_ dig_ctrl_inst.latch_mem_inst.RAM\[53\]\[0\]
+ _0154_ _0335_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_0_333 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[23\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND net179 dig_ctrl_inst.latch_mem_inst.gclk\[23\] dig_ctrl_inst.latch_mem_inst.RAM\[23\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
X_2224_ VGND VDPWR VDPWR VGND net160 _0868_ _0850_ sky130_fd_sc_hd__or2_1
X_2155_ VGND VDPWR VDPWR VGND _0775_ _0801_ _0782_ _0796_ net161 _0800_ sky130_fd_sc_hd__o221a_1
X_2086_ VDPWR VGND VDPWR VGND _0739_ _0732_ _0744_ _0737_ _0743_ sky130_fd_sc_hd__or4_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[12\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND net196 dig_ctrl_inst.latch_mem_inst.gclk\[12\] dig_ctrl_inst.latch_mem_inst.RAM\[12\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
X_1939_ VDPWR VGND VDPWR VGND net81 _0599_ dig_ctrl_inst.latch_mem_inst.RAM\[58\]\[5\]
+ net43 sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[5\].gen_latches\[7\].p_latch VGND VDPWR VDPWR
+ VGND net182 dig_ctrl_inst.latch_mem_inst.gclk\[5\] dig_ctrl_inst.latch_mem_inst.RAM\[5\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[39\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND net232 dig_ctrl_inst.latch_mem_inst.gclk\[39\] dig_ctrl_inst.latch_mem_inst.RAM\[39\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_11_Right_11 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.genblk1\[48\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[48\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[48\]._gclk clknet_leaf_13_clk sky130_fd_sc_hd__dlclkp_1
XPHY_EDGE_ROW_20_Right_20 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_1_119 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_1724_ VGND VDPWR VDPWR VGND _0385_ _0388_ _0387_ dig_ctrl_inst.latch_mem_inst.RAM\[23\]\[1\]
+ _0128_ _0386_ sky130_fd_sc_hd__a2111o_1
X_1655_ VGND VDPWR VDPWR VGND _0317_ _0320_ _0319_ dig_ctrl_inst.latch_mem_inst.RAM\[63\]\[0\]
+ _0163_ _0318_ sky130_fd_sc_hd__a2111o_1
X_1586_ VGND VDPWR VDPWR VGND _0252_ _1162_ net158 sky130_fd_sc_hd__nand2b_1
XFILLER_0_0_141 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
Xdig_ctrl_inst.latch_mem_inst.gen_words\[16\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND net189 dig_ctrl_inst.latch_mem_inst.gclk\[16\] dig_ctrl_inst.latch_mem_inst.RAM\[16\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
X_2069_ VDPWR VGND VDPWR VGND net111 _0727_ dig_ctrl_inst.latch_mem_inst.RAM\[34\]\[7\]
+ net49 sky130_fd_sc_hd__and3_2
X_2138_ VGND VDPWR VDPWR VGND _0784_ _0783_ net149 sky130_fd_sc_hd__nand2_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[50\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[50\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[50\]._gclk clknet_leaf_13_clk sky130_fd_sc_hd__dlclkp_1
X_2207_ VGND VDPWR VDPWR VGND _0851_ _0764_ _0815_ _0852_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_280 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
Xdig_ctrl_inst.latch_mem_inst.genblk1\[24\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[24\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[24\]._gclk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_54_169 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1440_ VDPWR VGND VDPWR VGND net107 _0153_ net137 net46 sky130_fd_sc_hd__and3_2
XFILLER_0_49_47 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1371_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[15\] _0119_ net143
+ sky130_fd_sc_hd__and2_1
XFILLER_0_77_228 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_45_169 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_136 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
X_1707_ VGND VDPWR VDPWR VGND _0371_ net106 dig_ctrl_inst.latch_mem_inst.RAM\[7\]\[1\]
+ net128 net102 sky130_fd_sc_hd__and4_1
X_1638_ VDPWR VGND VDPWR VGND net126 _0303_ dig_ctrl_inst.latch_mem_inst.RAM\[4\]\[0\]
+ net97 sky130_fd_sc_hd__and3_2
XPHY_EDGE_ROW_18_Left_96 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1569_ VGND VDPWR VDPWR VGND net158 _0235_ _1162_ sky130_fd_sc_hd__nor2_1
Xfanout98 VGND VDPWR VDPWR VGND net99 net98 sky130_fd_sc_hd__clkbuf_2
Xfanout65 VDPWR VGND VDPWR VGND net65 net70 sky130_fd_sc_hd__buf_2
Xfanout54 VGND VDPWR VDPWR VGND _0134_ net54 sky130_fd_sc_hd__clkbuf_2
Xfanout43 VGND VDPWR VDPWR VGND net44 net43 sky130_fd_sc_hd__clkbuf_2
Xfanout76 VDPWR VGND VDPWR VGND net76 net80 sky130_fd_sc_hd__buf_2
Xfanout87 VDPWR VGND VDPWR VGND net87 _1186_ sky130_fd_sc_hd__buf_2
XFILLER_0_36_136 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2472_ VGND VDPWR VDPWR VGND dig_ctrl_inst.synchronizer_port_i_inst\[1\].pipe\[0\]
+ net169 net4 clknet_leaf_5_clk sky130_fd_sc_hd__dfrtp_1
Xclkload13 VDPWR VGND VDPWR VGND clknet_leaf_6_clk clkload13/Y sky130_fd_sc_hd__clkinvlp_4
X_2610_ VGND VDPWR VDPWR VGND net24 dig_ctrl_inst.spi_miso_o sky130_fd_sc_hd__clkbuf_1
X_2541_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[2\]\[5\] net156 _0067_
+ clknet_leaf_7_clk sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_191 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_1354_ VDPWR VGND VDPWR VGND net145 dig_ctrl_inst.latch_mem_inst.data_we\[8\] net130
+ net86 sky130_fd_sc_hd__and3_2
X_1423_ VDPWR VGND VDPWR VGND _0145_ net53 net82 sky130_fd_sc_hd__and2_1
X_1285_ VGND VDPWR VDPWR VGND net250 dig_ctrl_inst.cpu_inst.regs\[1\]\[2\] _1127_
+ net254 sky130_fd_sc_hd__and3b_1
XFILLER_0_41_92 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xclkload7 VGND VDPWR VDPWR VGND clkload7/Y clknet_leaf_17_clk sky130_fd_sc_hd__inv_16
XFILLER_0_18_125 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xfanout222 VDPWR VGND VDPWR VGND net222 net227 sky130_fd_sc_hd__buf_2
Xfanout200 VGND VDPWR VDPWR VGND net201 net200 sky130_fd_sc_hd__clkbuf_2
Xfanout211 VDPWR VGND VDPWR VGND net211 net214 sky130_fd_sc_hd__buf_2
Xfanout233 VGND VDPWR VDPWR VGND net234 net233 sky130_fd_sc_hd__clkbuf_2
Xfanout266 VGND VDPWR VDPWR VGND net266 net14 sky130_fd_sc_hd__buf_1
Xfanout244 VGND VDPWR VDPWR VGND net286 net244 sky130_fd_sc_hd__clkbuf_2
Xfanout255 VGND VDPWR VDPWR VGND net256 net255 sky130_fd_sc_hd__clkbuf_2
X_1972_ VGND VDPWR VDPWR VGND _0596_ _0632_ _0613_ dig_ctrl_inst.latch_mem_inst.RAM\[7\]\[5\]
+ _1184_ _0611_ sky130_fd_sc_hd__a2111o_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[4\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[4\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[4\]._gclk sky130_fd_sc_hd__clkbuf_4
X_2455_ VGND VDPWR VDPWR VGND net335 _1032_ _1034_ _0112_ sky130_fd_sc_hd__mux2_1
X_2524_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[0\]\[4\] net157 _0050_
+ clknet_leaf_7_clk sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_49_Right_49 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_23_183 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
Xdig_ctrl_inst.latch_mem_inst.gen_words\[53\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND net181 dig_ctrl_inst.latch_mem_inst.gclk\[53\] dig_ctrl_inst.latch_mem_inst.RAM\[53\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
X_1406_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[33\] _0136_ net147
+ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_58_Right_58 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2386_ VGND VDPWR VDPWR VGND _1003_ _0997_ net315 _0074_ sky130_fd_sc_hd__mux2_1
Xhold19 VGND VDPWR VDPWR VGND dig_ctrl_inst.synchronizer_port_i_inst\[5\].pipe\[0\]
+ net301 sky130_fd_sc_hd__dlygate4sd3_1
X_1337_ VDPWR VGND VDPWR VGND _1177_ _1139_ _1123_ _1106_ _1090_ _1052_ sky130_fd_sc_hd__o2111a_1
X_1268_ VGND VDPWR VDPWR VGND _1110_ net250 dig_ctrl_inst.cpu_inst.regs\[1\]\[3\]
+ sky130_fd_sc_hd__nand2b_1
X_1199_ VDPWR VGND VDPWR VGND dig_ctrl_inst.spi_addr\[2\] _1043_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_67_Right_67 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[42\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND net199 dig_ctrl_inst.latch_mem_inst.gclk\[42\] dig_ctrl_inst.latch_mem_inst.RAM\[42\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_76_Right_76 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.genblk1\[17\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[17\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[17\]._gclk sky130_fd_sc_hd__clkbuf_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[31\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND net213 dig_ctrl_inst.latch_mem_inst.gclk\[31\] dig_ctrl_inst.latch_mem_inst.RAM\[31\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[20\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND net233 dig_ctrl_inst.latch_mem_inst.gclk\[20\] dig_ctrl_inst.latch_mem_inst.RAM\[20\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_4_309 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_37_231 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_2171_ VDPWR VGND VDPWR VGND net247 _0817_ net246 _0804_ sky130_fd_sc_hd__and3_2
X_2240_ VGND VDPWR VDPWR VGND net150 _0799_ _0798_ _0883_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_337 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_73_57 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
Xdig_ctrl_inst.latch_mem_inst.genblk1\[55\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[55\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[55\]._gclk clknet_leaf_19_clk sky130_fd_sc_hd__dlclkp_1
X_1886_ VGND VDPWR VDPWR VGND _0528_ _0547_ _0537_ dig_ctrl_inst.latch_mem_inst.RAM\[49\]\[4\]
+ _0152_ _0535_ sky130_fd_sc_hd__a2111o_1
X_1955_ VGND VDPWR VDPWR VGND _0615_ net116 dig_ctrl_inst.latch_mem_inst.RAM\[9\]\[5\]
+ net124 net88 sky130_fd_sc_hd__and4_1
XFILLER_0_3_331 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_28_297 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2438_ VGND VDPWR VDPWR VGND dig_ctrl_inst.mode_sync net171 dig_ctrl_inst.spi_receiver_inst.stb_o
+ _1048_ _1023_ sky130_fd_sc_hd__o211a_1
X_2507_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.instr\[6\] net151 _0033_ clknet_leaf_13_clk
+ sky130_fd_sc_hd__dfrtp_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[2\].gen_latches\[1\].p_latch VGND VDPWR VDPWR
+ VGND net229 dig_ctrl_inst.latch_mem_inst.gclk\[2\] dig_ctrl_inst.latch_mem_inst.RAM\[2\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
X_2369_ VGND VDPWR VDPWR VGND _0988_ _1000_ _0766_ sky130_fd_sc_hd__nor2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[46\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND net191 dig_ctrl_inst.latch_mem_inst.gclk\[46\] dig_ctrl_inst.latch_mem_inst.RAM\[46\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[35\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND net205 dig_ctrl_inst.latch_mem_inst.gclk\[35\] dig_ctrl_inst.latch_mem_inst.RAM\[35\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[24\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND net226 dig_ctrl_inst.latch_mem_inst.gclk\[24\] dig_ctrl_inst.latch_mem_inst.RAM\[24\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_57_337 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_6_Left_84 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1671_ VDPWR VGND VDPWR VGND net96 _0336_ dig_ctrl_inst.latch_mem_inst.RAM\[54\]\[0\]
+ net41 sky130_fd_sc_hd__and3_2
X_1740_ VGND VDPWR VDPWR VGND _0400_ _0403_ _0402_ dig_ctrl_inst.latch_mem_inst.RAM\[55\]\[2\]
+ _0155_ _0401_ sky130_fd_sc_hd__a2111o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[13\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND net240 dig_ctrl_inst.latch_mem_inst.gclk\[13\] dig_ctrl_inst.latch_mem_inst.RAM\[13\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
X_2085_ VDPWR VGND VDPWR VGND _0741_ _0728_ _0743_ _0740_ _0742_ sky130_fd_sc_hd__or4_1
X_2223_ VGND VDPWR VDPWR VGND _0247_ _0818_ _0867_ _0866_ _0864_ sky130_fd_sc_hd__o211ai_1
X_2154_ VGND VDPWR VDPWR VGND net149 _0799_ _0798_ _0800_ sky130_fd_sc_hd__mux2_1
X_1869_ VDPWR VGND VDPWR VGND net73 _0530_ dig_ctrl_inst.latch_mem_inst.RAM\[60\]\[4\]
+ net45 sky130_fd_sc_hd__and3_2
X_1938_ VDPWR VGND VDPWR VGND net111 _0598_ dig_ctrl_inst.latch_mem_inst.RAM\[34\]\[5\]
+ net48 sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[6\].gen_latches\[2\].p_latch VGND VDPWR VDPWR
+ VGND net222 dig_ctrl_inst.latch_mem_inst.gclk\[6\] dig_ctrl_inst.latch_mem_inst.RAM\[6\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_39_337 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_66_123 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[39\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND net199 dig_ctrl_inst.latch_mem_inst.gclk\[39\] dig_ctrl_inst.latch_mem_inst.RAM\[39\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[28\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND net216 dig_ctrl_inst.latch_mem_inst.gclk\[28\] dig_ctrl_inst.latch_mem_inst.RAM\[28\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[17\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND net233 dig_ctrl_inst.latch_mem_inst.gclk\[17\] dig_ctrl_inst.latch_mem_inst.RAM\[17\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
X_1723_ VGND VDPWR VDPWR VGND _0387_ net91 dig_ctrl_inst.latch_mem_inst.RAM\[59\]\[1\]
+ net106 net44 sky130_fd_sc_hd__and4_1
X_1654_ VDPWR VGND VDPWR VGND net128 _0319_ dig_ctrl_inst.latch_mem_inst.RAM\[6\]\[0\]
+ net94 sky130_fd_sc_hd__and3_2
X_2206_ VGND VDPWR VDPWR VGND _0851_ _0850_ _0849_ sky130_fd_sc_hd__nand2_1
X_1585_ VGND VDPWR VDPWR VGND _1147_ _0251_ _1153_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_153 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_131 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_2068_ VDPWR VGND VDPWR VGND net133 _0726_ dig_ctrl_inst.latch_mem_inst.RAM\[48\]\[7\]
+ net38 sky130_fd_sc_hd__and3_2
X_2137_ VGND VDPWR VDPWR VGND _0783_ _0777_ _0227_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_292 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
Xdig_ctrl_inst.latch_mem_inst.genblk1\[63\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[63\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[63\]._gclk sky130_fd_sc_hd__clkbuf_4
X_1370_ VGND VDPWR VDPWR VGND net128 net110 net77 _0119_ sky130_fd_sc_hd__and3_4
X_1706_ VGND VDPWR VDPWR VGND _0370_ net114 dig_ctrl_inst.latch_mem_inst.RAM\[14\]\[1\]
+ net128 net77 sky130_fd_sc_hd__and4_1
X_1637_ VGND VDPWR VDPWR VGND _0302_ net104 dig_ctrl_inst.latch_mem_inst.RAM\[35\]\[0\]
+ net138 net52 sky130_fd_sc_hd__and4_1
X_1499_ VDPWR VGND VDPWR VGND _1066_ _1062_ _0187_ _1064_ _0186_ sky130_fd_sc_hd__or4_2
X_1568_ VGND VDPWR VDPWR VGND _0234_ net158 _1162_ sky130_fd_sc_hd__nand2_1
Xfanout44 VDPWR VGND VDPWR VGND net44 _0150_ sky130_fd_sc_hd__buf_2
Xfanout55 VGND VDPWR VDPWR VGND net58 net55 sky130_fd_sc_hd__clkbuf_2
Xfanout99 VGND VDPWR VDPWR VGND net100 net99 sky130_fd_sc_hd__clkbuf_2
Xfanout77 VDPWR VGND VDPWR VGND net77 net80 sky130_fd_sc_hd__buf_2
Xfanout66 VGND VDPWR VDPWR VGND net69 net66 sky130_fd_sc_hd__clkbuf_2
Xfanout88 VDPWR VGND VDPWR VGND net88 net92 sky130_fd_sc_hd__buf_2
XFILLER_0_3_3 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
Xdig_ctrl_inst.latch_mem_inst.gen_words\[61\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND net215 dig_ctrl_inst.latch_mem_inst.gclk\[61\] dig_ctrl_inst.latch_mem_inst.RAM\[61\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
X_2471_ VGND VDPWR VDPWR VGND dig_ctrl_inst.synchronizer_port_i_inst\[2\].out net169
+ net303 clknet_leaf_4_clk sky130_fd_sc_hd__dfrtp_1
X_2540_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[2\]\[4\] net157 _0066_
+ clknet_leaf_6_clk sky130_fd_sc_hd__dfrtp_1
Xclkload14 VGND VDPWR VDPWR VGND clkload14/Y clknet_leaf_7_clk sky130_fd_sc_hd__clkinv_16
X_1422_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[41\] _0144_ net142
+ sky130_fd_sc_hd__and2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[50\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND net230 dig_ctrl_inst.latch_mem_inst.gclk\[50\] dig_ctrl_inst.latch_mem_inst.RAM\[50\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
X_1353_ VDPWR VGND VDPWR VGND net132 _1187_ net84 sky130_fd_sc_hd__and2_2
X_1284_ VGND VDPWR VDPWR VGND net254 net250 _1126_ dig_ctrl_inst.cpu_inst.regs\[2\]\[2\]
+ sky130_fd_sc_hd__and3b_1
Xclkload8 VGND VDPWR VDPWR VGND clknet_leaf_0_clk clkload8/Y sky130_fd_sc_hd__inv_8
Xdig_ctrl_inst.latch_mem_inst.genblk1\[62\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[62\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[62\]._gclk clknet_leaf_16_clk sky130_fd_sc_hd__dlclkp_1
Xfanout245 VDPWR VGND VDPWR VGND net245 dig_ctrl_inst.cpu_inst.cpu_state\[2\] sky130_fd_sc_hd__buf_2
Xfanout201 VDPWR VGND VDPWR VGND net201 net202 sky130_fd_sc_hd__buf_2
Xfanout234 VGND VDPWR VDPWR VGND net235 net234 sky130_fd_sc_hd__clkbuf_2
Xfanout223 VGND VDPWR VDPWR VGND net227 net223 sky130_fd_sc_hd__clkbuf_2
Xfanout212 VGND VDPWR VDPWR VGND net213 net212 sky130_fd_sc_hd__clkbuf_2
Xfanout256 VDPWR VGND VDPWR VGND dig_ctrl_inst.cpu_inst.arg1\[0\] net256 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_49_295 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1971_ VDPWR VGND VDPWR VGND _0629_ _0626_ _0631_ _0628_ _0630_ sky130_fd_sc_hd__or4_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[54\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND net219 dig_ctrl_inst.latch_mem_inst.gclk\[54\] dig_ctrl_inst.latch_mem_inst.RAM\[54\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
X_1405_ VGND VDPWR VDPWR VGND net136 net121 net56 _0136_ sky130_fd_sc_hd__and3_4
X_2454_ VGND VDPWR VDPWR VGND _1034_ _1025_ dig_ctrl_inst.spi_addr\[3\] dig_ctrl_inst.spi_addr\[4\]
+ _1027_ sky130_fd_sc_hd__and4_1
XFILLER_0_23_173 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2523_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[0\]\[3\] net154 _0049_
+ clknet_leaf_11_clk sky130_fd_sc_hd__dfrtp_2
X_2385_ VGND VDPWR VDPWR VGND _1003_ _0996_ net353 _0073_ sky130_fd_sc_hd__mux2_1
X_1336_ VGND VDPWR VDPWR VGND _1176_ _1052_ _1106_ _1090_ sky130_fd_sc_hd__o21a_1
X_1198_ VDPWR VGND VDPWR VGND net346 _1042_ sky130_fd_sc_hd__inv_2
Xinput1 VGND VDPWR VDPWR VGND net1 port_ms_i sky130_fd_sc_hd__buf_1
X_1267_ VGND VDPWR VDPWR VGND net254 _1109_ net250 dig_ctrl_inst.cpu_inst.regs\[3\]\[3\]
+ sky130_fd_sc_hd__nand3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[43\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND net239 dig_ctrl_inst.latch_mem_inst.gclk\[43\] dig_ctrl_inst.latch_mem_inst.RAM\[43\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[56\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[56\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[56\]._gclk sky130_fd_sc_hd__clkbuf_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[31\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND net185 dig_ctrl_inst.latch_mem_inst.gclk\[31\] dig_ctrl_inst.latch_mem_inst.RAM\[31\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_32_29 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_37_243 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
Xdig_ctrl_inst.latch_mem_inst.gen_words\[20\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND net199 dig_ctrl_inst.latch_mem_inst.gclk\[20\] dig_ctrl_inst.latch_mem_inst.RAM\[20\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_20_132 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_73_69 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
X_2170_ VGND VDPWR VDPWR VGND net165 _0815_ _0764_ _0816_ sky130_fd_sc_hd__mux2_1
X_1954_ VDPWR VGND VDPWR VGND net113 _0614_ dig_ctrl_inst.latch_mem_inst.RAM\[50\]\[5\]
+ net46 sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[58\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND net214 dig_ctrl_inst.latch_mem_inst.gclk\[58\] dig_ctrl_inst.latch_mem_inst.RAM\[58\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_43_202 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1885_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[11\]\[4\] _0113_ _0546_
+ dig_ctrl_inst.latch_mem_inst.RAM\[39\]\[4\] _0142_ sky130_fd_sc_hd__a22o_1
X_2368_ VGND VDPWR VDPWR VGND _0991_ _0999_ dig_ctrl_inst.cpu_inst.regs\[1\]\[6\]
+ _0060_ sky130_fd_sc_hd__mux2_1
X_2437_ VDPWR VGND VDPWR VGND _1022_ _1048_ dig_ctrl_inst.mode_sync sky130_fd_sc_hd__and2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[47\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND net232 dig_ctrl_inst.latch_mem_inst.gclk\[47\] dig_ctrl_inst.latch_mem_inst.RAM\[47\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_44_3 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_2506_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.instr\[5\] net151 _0032_ clknet_leaf_13_clk
+ sky130_fd_sc_hd__dfrtp_1
X_1319_ VDPWR VGND VDPWR VGND net256 _1161_ net252 dig_ctrl_inst.cpu_inst.regs\[0\]\[4\]
+ sky130_fd_sc_hd__or3_1
X_2299_ VDPWR VGND VDPWR VGND _0940_ _0812_ _1147_ _0227_ _0807_ _0939_ sky130_fd_sc_hd__a221o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[2\].gen_latches\[5\].p_latch VGND VDPWR VDPWR
+ VGND net195 dig_ctrl_inst.latch_mem_inst.gclk\[2\] dig_ctrl_inst.latch_mem_inst.RAM\[2\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_68_25 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1670_ VGND VDPWR VDPWR VGND _0335_ net117 dig_ctrl_inst.latch_mem_inst.RAM\[9\]\[0\]
+ net125 net89 sky130_fd_sc_hd__and4_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[24\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND net186 dig_ctrl_inst.latch_mem_inst.gclk\[24\] dig_ctrl_inst.latch_mem_inst.RAM\[24\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
X_2222_ VDPWR VGND VDPWR VGND dig_ctrl_inst.cpu_inst.data\[2\] _0865_ _0866_ _0813_
+ sky130_fd_sc_hd__a21oi_1
X_2084_ VGND VDPWR VDPWR VGND _0718_ _0742_ _0729_ dig_ctrl_inst.latch_mem_inst.RAM\[17\]\[7\]
+ _0122_ _0721_ sky130_fd_sc_hd__a2111o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[13\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND net203 dig_ctrl_inst.latch_mem_inst.gclk\[13\] dig_ctrl_inst.latch_mem_inst.RAM\[13\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
X_2153_ VGND VDPWR VDPWR VGND _0799_ net140 net160 sky130_fd_sc_hd__nand2_1
X_1937_ VDPWR VGND VDPWR VGND net99 _0597_ dig_ctrl_inst.latch_mem_inst.RAM\[20\]\[5\]
+ net66 sky130_fd_sc_hd__and3_2
X_1799_ VDPWR VGND VDPWR VGND _0428_ _0462_ _0461_ _0279_ dig_ctrl_inst.latch_mem_inst.RAM\[0\]\[2\]
+ sky130_fd_sc_hd__o2bb2a_1
X_1868_ VGND VDPWR VDPWR VGND _0529_ net75 dig_ctrl_inst.latch_mem_inst.RAM\[63\]\[4\]
+ net104 net39 sky130_fd_sc_hd__and4_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[6\].gen_latches\[6\].p_latch VGND VDPWR VDPWR
+ VGND net194 dig_ctrl_inst.latch_mem_inst.gclk\[6\] dig_ctrl_inst.latch_mem_inst.RAM\[6\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[28\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND net181 dig_ctrl_inst.latch_mem_inst.gclk\[28\] dig_ctrl_inst.latch_mem_inst.RAM\[28\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
X_1722_ VDPWR VGND VDPWR VGND net135 _0386_ dig_ctrl_inst.latch_mem_inst.RAM\[48\]\[1\]
+ net44 sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[17\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND net200 dig_ctrl_inst.latch_mem_inst.gclk\[17\] dig_ctrl_inst.latch_mem_inst.RAM\[17\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
X_1653_ VGND VDPWR VDPWR VGND _0318_ net114 dig_ctrl_inst.latch_mem_inst.RAM\[14\]\[0\]
+ net128 net75 sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_9_Right_9 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1584_ VDPWR VGND VDPWR VGND _0249_ _0237_ _0236_ _0250_ sky130_fd_sc_hd__a21o_1
XFILLER_0_28_61 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_2205_ VGND VDPWR VDPWR VGND net165 _0850_ net164 sky130_fd_sc_hd__or2_1
XFILLER_0_0_165 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.genblk1\[49\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[49\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[49\]._gclk sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_22_Left_100 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2067_ VDPWR VGND VDPWR VGND net124 _0725_ dig_ctrl_inst.latch_mem_inst.RAM\[10\]\[7\]
+ net83 sky130_fd_sc_hd__and3_2
X_2136_ VDPWR VGND VDPWR VGND _0775_ _0782_ _1099_ sky130_fd_sc_hd__or2_2
XFILLER_0_8_276 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_2604__270 VGND VDPWR VDPWR VGND net270 _2604__270/HI sky130_fd_sc_hd__conb_1
XFILLER_0_24_19 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_2611__274 VGND VDPWR VDPWR VGND net274 _2611__274/HI sky130_fd_sc_hd__conb_1
XFILLER_0_54_149 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_62_193 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_49_38 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_4_29 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1705_ VGND VDPWR VDPWR VGND _0366_ _0369_ _0368_ dig_ctrl_inst.latch_mem_inst.RAM\[51\]\[1\]
+ _0153_ _0367_ sky130_fd_sc_hd__a2111o_1
X_1636_ VGND VDPWR VDPWR VGND _0301_ net103 dig_ctrl_inst.latch_mem_inst.RAM\[23\]\[0\]
+ net104 net62 sky130_fd_sc_hd__and4_1
X_1567_ VDPWR VGND VDPWR VGND _0233_ net158 _1162_ sky130_fd_sc_hd__and2_1
X_1498_ VDPWR VGND VDPWR VGND _1036_ _0186_ _1037_ net245 sky130_fd_sc_hd__or3_4
X_2119_ VDPWR VGND VDPWR VGND net248 _0765_ dig_ctrl_inst.cpu_inst.instr\[6\] dig_ctrl_inst.cpu_inst.instr\[7\]
+ sky130_fd_sc_hd__or3_1
Xfanout56 VGND VDPWR VDPWR VGND net57 net56 sky130_fd_sc_hd__clkbuf_2
Xfanout45 VDPWR VGND VDPWR VGND net45 net47 sky130_fd_sc_hd__buf_2
Xfanout67 VGND VDPWR VDPWR VGND net69 net67 sky130_fd_sc_hd__clkbuf_2
Xfanout78 VGND VDPWR VDPWR VGND net80 net78 sky130_fd_sc_hd__clkbuf_2
Xfanout89 VGND VDPWR VDPWR VGND net92 net89 sky130_fd_sc_hd__clkbuf_2
Xclkload15 VGND VDPWR VDPWR VGND clkload15/Y clknet_leaf_8_clk sky130_fd_sc_hd__inv_16
Xdig_ctrl_inst.latch_mem_inst.gen_words\[61\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND net184 dig_ctrl_inst.latch_mem_inst.gclk\[61\] dig_ctrl_inst.latch_mem_inst.RAM\[61\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[20\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[20\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[20\]._gclk sky130_fd_sc_hd__clkbuf_4
X_2470_ VGND VDPWR VDPWR VGND dig_ctrl_inst.synchronizer_port_i_inst\[2\].pipe\[0\]
+ net169 net5 clknet_leaf_5_clk sky130_fd_sc_hd__dfrtp_1
X_1421_ VDPWR VGND VDPWR VGND net88 _0144_ net116 net49 sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[50\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND net202 dig_ctrl_inst.latch_mem_inst.gclk\[50\] dig_ctrl_inst.latch_mem_inst.RAM\[50\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
X_1352_ VDPWR VGND VDPWR VGND _1186_ _1139_ _1122_ _1107_ _1090_ _1052_ sky130_fd_sc_hd__o2111a_1
X_1283_ VDPWR VGND VDPWR VGND net250 _1125_ net254 dig_ctrl_inst.cpu_inst.regs\[3\]\[2\]
+ sky130_fd_sc_hd__and3_2
Xclkload9 VGND VDPWR VDPWR VGND clknet_leaf_1_clk clkload9/Y sky130_fd_sc_hd__inv_12
Xfanout202 VDPWR VGND VDPWR VGND net202 net287 sky130_fd_sc_hd__buf_2
Xfanout235 VDPWR VGND VDPWR VGND net290 net235 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout224 VGND VDPWR VDPWR VGND net226 net224 sky130_fd_sc_hd__clkbuf_2
X_1619_ VGND VDPWR VDPWR VGND _0284_ net79 dig_ctrl_inst.latch_mem_inst.RAM\[47\]\[0\]
+ net106 net53 sky130_fd_sc_hd__and4_1
XFILLER_0_1_293 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
Xfanout246 VDPWR VGND VDPWR VGND net246 dig_ctrl_inst.cpu_inst.instr\[5\] sky130_fd_sc_hd__buf_2
Xfanout213 VDPWR VGND VDPWR VGND net213 net214 sky130_fd_sc_hd__buf_2
Xfanout257 VGND VDPWR VDPWR VGND net260 net257 sky130_fd_sc_hd__clkbuf_2
X_2599_ VDPWR VGND VDPWR VGND net15 clknet_leaf_12_clk sky130_fd_sc_hd__buf_2
XFILLER_0_66_91 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_1970_ VGND VDPWR VDPWR VGND _0588_ _0630_ _0617_ dig_ctrl_inst.latch_mem_inst.RAM\[5\]\[5\]
+ _0272_ _0591_ sky130_fd_sc_hd__a2111o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[54\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND net188 dig_ctrl_inst.latch_mem_inst.gclk\[54\] dig_ctrl_inst.latch_mem_inst.RAM\[54\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
X_2522_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[0\]\[2\] net154 _0048_
+ clknet_leaf_11_clk sky130_fd_sc_hd__dfrtp_1
X_1335_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[1\] _1175_ net144
+ sky130_fd_sc_hd__and2_1
X_2453_ VDPWR VGND VDPWR VGND _0111_ _1033_ _1032_ sky130_fd_sc_hd__and2_1
X_1404_ VDPWR VGND VDPWR VGND net143 dig_ctrl_inst.latch_mem_inst.data_we\[32\] net134
+ net50 sky130_fd_sc_hd__and3_2
X_2384_ VGND VDPWR VDPWR VGND _1003_ _0995_ net319 _0072_ sky130_fd_sc_hd__mux2_1
Xinput2 VGND VDPWR VDPWR VGND net2 rst_n sky130_fd_sc_hd__clkbuf_1
X_1197_ VDPWR VGND VDPWR VGND net264 _1041_ sky130_fd_sc_hd__inv_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[43\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND net205 dig_ctrl_inst.latch_mem_inst.gclk\[43\] dig_ctrl_inst.latch_mem_inst.RAM\[43\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
X_1266_ VGND VDPWR VDPWR VGND _1108_ _1070_ _1072_ _1054_ _1045_ sky130_fd_sc_hd__a211o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[32\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND net220 dig_ctrl_inst.latch_mem_inst.gclk\[32\] dig_ctrl_inst.latch_mem_inst.RAM\[32\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[21\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND net240 dig_ctrl_inst.latch_mem_inst.gclk\[21\] dig_ctrl_inst.latch_mem_inst.RAM\[21\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_37_255 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_20_144 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_69_Left_147 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_43_214 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
Xdig_ctrl_inst.latch_mem_inst.gen_words\[58\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND net183 dig_ctrl_inst.latch_mem_inst.gclk\[58\] dig_ctrl_inst.latch_mem_inst.RAM\[58\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
X_1953_ VGND VDPWR VDPWR VGND _0613_ net90 dig_ctrl_inst.latch_mem_inst.RAM\[27\]\[5\]
+ net107 net68 sky130_fd_sc_hd__and4_1
X_1884_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[22\]\[4\] _0127_ _0545_
+ dig_ctrl_inst.latch_mem_inst.RAM\[53\]\[4\] _0154_ sky130_fd_sc_hd__a22o_1
X_2505_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.instr\[4\] net151 _0031_ clknet_leaf_14_clk
+ sky130_fd_sc_hd__dfrtp_1
X_2436_ VGND VDPWR VDPWR VGND _0106_ _1015_ _0195_ _1020_ sky130_fd_sc_hd__o21a_1
X_1318_ VGND VDPWR VDPWR VGND _1160_ net252 dig_ctrl_inst.cpu_inst.regs\[1\]\[4\]
+ sky130_fd_sc_hd__and2b_1
X_2367_ VDPWR VGND VDPWR VGND _0766_ _0999_ _0967_ _0970_ sky130_fd_sc_hd__o21bai_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[3\].gen_latches\[0\].p_latch VGND VDPWR VDPWR
+ VGND net243 dig_ctrl_inst.latch_mem_inst.gclk\[3\] dig_ctrl_inst.latch_mem_inst.RAM\[3\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[47\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND net199 dig_ctrl_inst.latch_mem_inst.gclk\[47\] dig_ctrl_inst.latch_mem_inst.RAM\[47\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_37_3 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_2298_ VGND VDPWR VDPWR VGND _0939_ _0844_ _0937_ net158 _0938_ sky130_fd_sc_hd__a211o_1
X_1249_ VGND VDPWR VDPWR VGND _1091_ _1042_ net14 sky130_fd_sc_hd__nand2_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[0\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[0\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[0\]._gclk sky130_fd_sc_hd__clkbuf_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[36\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND net217 dig_ctrl_inst.latch_mem_inst.gclk\[36\] dig_ctrl_inst.latch_mem_inst.RAM\[36\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_34_258 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
Xdig_ctrl_inst.latch_mem_inst.gen_words\[25\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND net235 dig_ctrl_inst.latch_mem_inst.gclk\[25\] dig_ctrl_inst.latch_mem_inst.RAM\[25\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_input_latches\[1\].n_latch VGND VDPWR VDPWR VGND
+ dig_ctrl_inst.data_out\[1\] clknet_leaf_3_clk dig_ctrl_inst.latch_mem_inst.wdata\[1\]
+ sky130_fd_sc_hd__dlxtn_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[13\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[13\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[13\]._gclk sky130_fd_sc_hd__clkbuf_4
X_2152_ VGND VDPWR VDPWR VGND _0798_ net140 net163 sky130_fd_sc_hd__nand2_1
X_2221_ VDPWR VGND VDPWR VGND net163 _0812_ _0865_ net164 _0844_ sky130_fd_sc_hd__a22o_1
X_2083_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[41\]\[7\] _0144_ _0741_
+ dig_ctrl_inst.latch_mem_inst.RAM\[47\]\[7\] _0149_ sky130_fd_sc_hd__a22o_1
X_1936_ VGND VDPWR VDPWR VGND _0596_ net78 dig_ctrl_inst.latch_mem_inst.RAM\[47\]\[5\]
+ net107 net56 sky130_fd_sc_hd__and4_1
X_1867_ VGND VDPWR VDPWR VGND _0528_ net79 dig_ctrl_inst.latch_mem_inst.RAM\[30\]\[4\]
+ net115 net64 sky130_fd_sc_hd__and4_1
X_1798_ VGND VDPWR VDPWR VGND _0460_ _0443_ _0277_ _0271_ _0461_ sky130_fd_sc_hd__o211a_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[7\].gen_latches\[1\].p_latch VGND VDPWR VDPWR
+ VGND net234 dig_ctrl_inst.latch_mem_inst.gclk\[7\] dig_ctrl_inst.latch_mem_inst.RAM\[7\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
X_2419_ VGND VDPWR VDPWR VGND net139 dig_ctrl_inst.cpu_inst.port_o\[1\] net17 _0097_
+ sky130_fd_sc_hd__mux2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[29\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND net224 dig_ctrl_inst.latch_mem_inst.gclk\[29\] dig_ctrl_inst.latch_mem_inst.RAM\[29\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[18\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND net236 dig_ctrl_inst.latch_mem_inst.gclk\[18\] dig_ctrl_inst.latch_mem_inst.RAM\[18\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
X_1721_ VGND VDPWR VDPWR VGND _0385_ net77 dig_ctrl_inst.latch_mem_inst.RAM\[61\]\[1\]
+ net122 net44 sky130_fd_sc_hd__and4_1
X_1652_ VDPWR VGND VDPWR VGND net113 _0317_ dig_ctrl_inst.latch_mem_inst.RAM\[34\]\[0\]
+ net54 sky130_fd_sc_hd__and3_2
X_1583_ VGND VDPWR VDPWR VGND _0249_ _0248_ _0241_ sky130_fd_sc_hd__nand2_1
X_2204_ VGND VDPWR VDPWR VGND _0849_ net164 net165 sky130_fd_sc_hd__nand2_1
X_2135_ VGND VDPWR VDPWR VGND net149 _0780_ _0778_ _0781_ sky130_fd_sc_hd__mux2_1
X_2066_ VDPWR VGND VDPWR VGND net127 _0724_ dig_ctrl_inst.latch_mem_inst.RAM\[8\]\[7\]
+ net86 sky130_fd_sc_hd__and3_2
XFILLER_0_36_309 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1919_ VGND VDPWR VDPWR VGND _0579_ net101 dig_ctrl_inst.latch_mem_inst.RAM\[39\]\[5\]
+ net109 net55 sky130_fd_sc_hd__and4_1
XFILLER_0_8_72 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_53 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_18_309 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_1704_ VGND VDPWR VDPWR VGND _0368_ net102 dig_ctrl_inst.latch_mem_inst.RAM\[37\]\[1\]
+ net119 net57 sky130_fd_sc_hd__and4_1
XFILLER_0_30_41 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1635_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[37\]\[0\] _0140_ _0300_
+ dig_ctrl_inst.latch_mem_inst.RAM\[58\]\[0\] _0158_ sky130_fd_sc_hd__a22o_1
X_1566_ VGND VDPWR VDPWR VGND _0232_ _1153_ _0224_ _1147_ _0231_ sky130_fd_sc_hd__a211o_1
X_1497_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.cpu_state\[1\] _0185_ net245
+ dig_ctrl_inst.cpu_inst.cpu_state\[0\] sky130_fd_sc_hd__and3b_2
X_2049_ VGND VDPWR VDPWR VGND net35 net36 _0277_ _0271_ _0708_ sky130_fd_sc_hd__o211a_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[13\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[13\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[13\]._gclk clknet_leaf_16_clk sky130_fd_sc_hd__dlclkp_1
X_2118_ VGND VDPWR VDPWR VGND _1062_ _0764_ _1057_ sky130_fd_sc_hd__nor2_2
Xfanout57 VGND VDPWR VDPWR VGND net58 net57 sky130_fd_sc_hd__clkbuf_2
Xfanout46 VGND VDPWR VDPWR VGND net47 net46 sky130_fd_sc_hd__clkbuf_2
Xfanout68 VGND VDPWR VDPWR VGND net69 net68 sky130_fd_sc_hd__clkbuf_2
Xfanout79 VDPWR VGND VDPWR VGND net79 net80 sky130_fd_sc_hd__buf_2
XFILLER_0_32_301 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
Xdig_ctrl_inst.latch_mem_inst.gen_words\[62\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND net222 dig_ctrl_inst.latch_mem_inst.gclk\[62\] dig_ctrl_inst.latch_mem_inst.RAM\[62\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
Xclkload16 VGND VDPWR VDPWR VGND clkload16/Y clknet_leaf_9_clk sky130_fd_sc_hd__inv_16
Xdig_ctrl_inst.latch_mem_inst.gen_words\[51\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND net243 dig_ctrl_inst.latch_mem_inst.gclk\[51\] dig_ctrl_inst.latch_mem_inst.RAM\[51\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_41_Left_119 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1351_ VGND VDPWR VDPWR VGND _1138_ _1185_ _1123_ sky130_fd_sc_hd__nor2_1
XFILLER_0_50_153 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1420_ VDPWR VGND VDPWR VGND net84 dig_ctrl_inst.latch_mem_inst.data_we\[40\] net142
+ net49 sky130_fd_sc_hd__and3_2
XPHY_EDGE_ROW_50_Left_128 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1282_ VGND VDPWR VDPWR VGND _1053_ _1073_ _1071_ dig_ctrl_inst.cpu_inst.ip\[2\]
+ _1124_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_25_85 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_33_109 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1618_ VDPWR VGND VDPWR VGND net127 _0283_ dig_ctrl_inst.latch_mem_inst.RAM\[12\]\[0\]
+ net73 sky130_fd_sc_hd__and3_2
XFILLER_0_26_161 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_14_334 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_1_261 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_2598_ VDPWR VGND VDPWR VGND dig_ctrl_inst.spi_addr\[5\] clknet_leaf_3_clk _0112_
+ sky130_fd_sc_hd__dfxtp_1
Xfanout258 VDPWR VGND VDPWR VGND net258 net260 sky130_fd_sc_hd__buf_2
Xfanout225 VGND VDPWR VDPWR VGND net225 net226 sky130_fd_sc_hd__buf_1
Xfanout236 VGND VDPWR VDPWR VGND net244 net236 sky130_fd_sc_hd__clkbuf_2
Xfanout203 VGND VDPWR VDPWR VGND net204 net203 sky130_fd_sc_hd__clkbuf_2
Xfanout247 VDPWR VGND VDPWR VGND net247 dig_ctrl_inst.cpu_inst.instr\[4\] sky130_fd_sc_hd__buf_2
X_1549_ VGND VDPWR VDPWR VGND _0191_ net159 dig_ctrl_inst.cpu_inst.data\[5\] _0216_
+ sky130_fd_sc_hd__mux2_1
Xfanout214 VDPWR VGND VDPWR VGND net289 net214 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_32_197 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
Xdig_ctrl_inst.latch_mem_inst.gen_words\[55\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND net228 dig_ctrl_inst.latch_mem_inst.gclk\[55\] dig_ctrl_inst.latch_mem_inst.RAM\[55\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_11_337 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2521_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[0\]\[1\] net152 _0047_
+ clknet_leaf_12_clk sky130_fd_sc_hd__dfrtp_1
X_2452_ VGND VDPWR VDPWR VGND _1023_ dig_ctrl_inst.spi_addr\[4\] dig_ctrl_inst.spi_addr\[3\]
+ _1027_ _1033_ sky130_fd_sc_hd__a31o_1
X_1265_ VGND VDPWR VDPWR VGND _1105_ _1092_ net265 _1107_ _1091_ sky130_fd_sc_hd__o31ai_4
XPHY_EDGE_ROW_18_Right_18 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1403_ VDPWR VGND VDPWR VGND _0135_ net50 net134 sky130_fd_sc_hd__and2_1
X_1334_ VGND VDPWR VDPWR VGND net138 net125 net117 _1175_ sky130_fd_sc_hd__and3_4
X_2383_ VGND VDPWR VDPWR VGND _1003_ _0994_ net318 _0071_ sky130_fd_sc_hd__mux2_1
Xinput3 VGND VDPWR VDPWR VGND net3 ui_in[0] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_50 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1196_ VDPWR VGND VDPWR VGND dig_ctrl_inst.cpu_inst.ip\[0\] _1040_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_27_Right_27 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_36_Right_36 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[32\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND net186 dig_ctrl_inst.latch_mem_inst.gclk\[32\] dig_ctrl_inst.latch_mem_inst.RAM\[32\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_45_Right_45 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[21\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND net208 dig_ctrl_inst.latch_mem_inst.gclk\[21\] dig_ctrl_inst.latch_mem_inst.RAM\[21\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_54_Right_54 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[59\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND net223 dig_ctrl_inst.latch_mem_inst.gclk\[59\] dig_ctrl_inst.latch_mem_inst.RAM\[59\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[10\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND net222 dig_ctrl_inst.latch_mem_inst.gclk\[10\] dig_ctrl_inst.latch_mem_inst.RAM\[10\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_63_Right_63 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_73_27 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1883_ VDPWR VGND VDPWR VGND _0544_ _0153_ dig_ctrl_inst.latch_mem_inst.RAM\[46\]\[4\]
+ dig_ctrl_inst.latch_mem_inst.RAM\[51\]\[4\] _0148_ _0530_ sky130_fd_sc_hd__a221o_1
X_1952_ VDPWR VGND VDPWR VGND net94 _0612_ dig_ctrl_inst.latch_mem_inst.RAM\[38\]\[5\]
+ net57 sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[48\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND net239 dig_ctrl_inst.latch_mem_inst.gclk\[48\] dig_ctrl_inst.latch_mem_inst.RAM\[48\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
X_2435_ VGND VDPWR VDPWR VGND _1015_ dig_ctrl_inst.cpu_inst.cpu_state\[1\] _1073_
+ _0105_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_72_Right_72 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_51_281 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2504_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.arg1\[1\] net152 _0030_ clknet_leaf_11_clk
+ sky130_fd_sc_hd__dfrtp_1
X_1248_ VDPWR VGND VDPWR VGND _1074_ _1089_ _1081_ _1075_ _1090_ sky130_fd_sc_hd__o211a_2
X_2366_ VGND VDPWR VDPWR VGND _0991_ _0998_ net316 _0059_ sky130_fd_sc_hd__mux2_1
X_1317_ VGND VDPWR VDPWR VGND net256 net252 _1159_ dig_ctrl_inst.cpu_inst.regs\[2\]\[4\]
+ sky130_fd_sc_hd__and3b_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[3\].gen_latches\[4\].p_latch VGND VDPWR VDPWR
+ VGND net210 dig_ctrl_inst.latch_mem_inst.gclk\[3\] dig_ctrl_inst.latch_mem_inst.RAM\[3\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
X_2297_ VDPWR VGND VDPWR VGND _0938_ net248 _0804_ _0929_ _0930_ _1039_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_66_318 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[36\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND net180 dig_ctrl_inst.latch_mem_inst.gclk\[36\] dig_ctrl_inst.latch_mem_inst.RAM\[36\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[52\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[52\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[52\]._gclk sky130_fd_sc_hd__clkbuf_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[25\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND net196 dig_ctrl_inst.latch_mem_inst.gclk\[25\] dig_ctrl_inst.latch_mem_inst.RAM\[25\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_input_latches\[5\].n_latch VGND VDPWR VDPWR VGND
+ dig_ctrl_inst.data_out\[5\] clknet_leaf_3_clk dig_ctrl_inst.latch_mem_inst.wdata\[5\]
+ sky130_fd_sc_hd__dlxtn_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[14\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND net215 dig_ctrl_inst.latch_mem_inst.gclk\[14\] dig_ctrl_inst.latch_mem_inst.RAM\[14\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_0_337 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2082_ VGND VDPWR VDPWR VGND _0713_ _0740_ _0722_ dig_ctrl_inst.latch_mem_inst.RAM\[3\]\[7\]
+ _1180_ _0717_ sky130_fd_sc_hd__a2111o_1
X_2151_ VGND VDPWR VDPWR VGND _0775_ _0797_ net161 sky130_fd_sc_hd__nor2_1
X_2220_ VGND VDPWR VDPWR VGND _0805_ _0864_ _0810_ _0863_ _0245_ _0244_ sky130_fd_sc_hd__o221a_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[18\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[18\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[18\]._gclk clknet_leaf_16_clk sky130_fd_sc_hd__dlclkp_1
X_1797_ VGND VDPWR VDPWR VGND _0459_ _0455_ _0460_ _0447_ _0451_ sky130_fd_sc_hd__nor4_1
X_1935_ VGND VDPWR VDPWR VGND _0595_ net102 dig_ctrl_inst.latch_mem_inst.RAM\[21\]\[5\]
+ net119 net63 sky130_fd_sc_hd__and4_1
X_1866_ VDPWR VGND VDPWR VGND net71 _0527_ dig_ctrl_inst.latch_mem_inst.RAM\[44\]\[4\]
+ net48 sky130_fd_sc_hd__and3_2
X_2418_ VGND VDPWR VDPWR VGND net139 dig_ctrl_inst.cpu_inst.port_o\[0\] net16 _0096_
+ sky130_fd_sc_hd__mux2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[7\].gen_latches\[5\].p_latch VGND VDPWR VDPWR
+ VGND net201 dig_ctrl_inst.latch_mem_inst.gclk\[7\] dig_ctrl_inst.latch_mem_inst.RAM\[7\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
X_2349_ VDPWR VGND VDPWR VGND _0968_ _0988_ _0221_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_0_Right_0 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.genblk1\[20\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[20\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[20\]._gclk clknet_leaf_4_clk sky130_fd_sc_hd__dlclkp_1
XFILLER_0_54_29 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[29\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND net188 dig_ctrl_inst.latch_mem_inst.gclk\[29\] dig_ctrl_inst.latch_mem_inst.RAM\[29\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
X_1720_ VGND VDPWR VDPWR VGND _0381_ _0384_ _0383_ dig_ctrl_inst.latch_mem_inst.RAM\[35\]\[1\]
+ _0138_ _0382_ sky130_fd_sc_hd__a2111o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[18\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND net210 dig_ctrl_inst.latch_mem_inst.gclk\[18\] dig_ctrl_inst.latch_mem_inst.RAM\[18\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
X_1651_ VDPWR VGND VDPWR VGND _0316_ _0132_ dig_ctrl_inst.latch_mem_inst.RAM\[19\]\[0\]
+ dig_ctrl_inst.latch_mem_inst.RAM\[30\]\[0\] _0124_ _0315_ sky130_fd_sc_hd__a221o_1
X_1582_ VGND VDPWR VDPWR VGND _0248_ _0247_ net161 net160 _0242_ _0243_ sky130_fd_sc_hd__a32o_1
XFILLER_0_28_85 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2065_ VDPWR VGND VDPWR VGND net81 _0723_ dig_ctrl_inst.latch_mem_inst.RAM\[42\]\[7\]
+ net53 sky130_fd_sc_hd__and3_2
X_2134_ VGND VDPWR VDPWR VGND _0780_ net140 net158 sky130_fd_sc_hd__nand2_1
X_2203_ VGND VDPWR VDPWR VGND _0848_ _0807_ _0845_ _1098_ _0847_ sky130_fd_sc_hd__a211o_1
XFILLER_0_71_140 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1849_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[13\]\[3\] _0117_ _0511_
+ dig_ctrl_inst.latch_mem_inst.RAM\[31\]\[3\] _0133_ sky130_fd_sc_hd__a22o_1
X_1918_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[0\]\[5\] _0578_ _0271_
+ _0277_ sky130_fd_sc_hd__or3_1
X_1634_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[32\]\[0\] _0135_ _0299_
+ dig_ctrl_inst.latch_mem_inst.RAM\[36\]\[0\] _0139_ sky130_fd_sc_hd__a22o_1
X_1703_ VGND VDPWR VDPWR VGND _0367_ net77 dig_ctrl_inst.latch_mem_inst.RAM\[46\]\[1\]
+ net115 net57 sky130_fd_sc_hd__and4_1
Xclkbuf_leaf_11_clk VGND VDPWR VDPWR VGND clknet_leaf_11_clk clknet_1_0__leaf_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_39_51 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1496_ VDPWR VGND VDPWR VGND _0183_ _0184_ sky130_fd_sc_hd__inv_2
X_1565_ VGND VDPWR VDPWR VGND _0230_ _0231_ _0228_ sky130_fd_sc_hd__nor2_1
X_2117_ VGND VDPWR VDPWR VGND _1051_ net310 net245 _0045_ sky130_fd_sc_hd__mux2_1
X_2048_ VGND VDPWR VDPWR VGND _0706_ _0702_ _0707_ _0694_ _0698_ sky130_fd_sc_hd__nor4_1
Xfanout69 VGND VDPWR VDPWR VGND net70 net69 sky130_fd_sc_hd__clkbuf_2
Xfanout47 VDPWR VGND VDPWR VGND net47 _0150_ sky130_fd_sc_hd__buf_2
XFILLER_0_44_184 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
Xfanout58 VGND VDPWR VDPWR VGND _0134_ net58 sky130_fd_sc_hd__clkbuf_2
Xdig_ctrl_inst.latch_mem_inst.genblk1\[45\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[45\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[45\]._gclk sky130_fd_sc_hd__clkbuf_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[62\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND net187 dig_ctrl_inst.latch_mem_inst.gclk\[62\] dig_ctrl_inst.latch_mem_inst.RAM\[62\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
Xclkload17 VGND VDPWR VDPWR VGND clkload17/Y clknet_leaf_18_clk sky130_fd_sc_hd__clkinv_16
Xdig_ctrl_inst.latch_mem_inst.gen_words\[51\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND net207 dig_ctrl_inst.latch_mem_inst.gclk\[51\] dig_ctrl_inst.latch_mem_inst.RAM\[51\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_35_184 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1281_ VGND VDPWR VDPWR VGND _1123_ _1121_ net264 _1044_ _1108_ _1115_ sky130_fd_sc_hd__a32o_1
X_1350_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[7\] _1184_ net147
+ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_0_clk VGND VDPWR VDPWR VGND clknet_leaf_0_clk clknet_1_1__leaf_clk sky130_fd_sc_hd__clkbuf_8
Xdig_ctrl_inst.latch_mem_inst.gen_words\[40\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND net223 dig_ctrl_inst.latch_mem_inst.gclk\[40\] dig_ctrl_inst.latch_mem_inst.RAM\[40\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
X_2597_ VDPWR VGND VDPWR VGND dig_ctrl_inst.spi_addr\[4\] clknet_leaf_3_clk _0111_
+ sky130_fd_sc_hd__dfxtp_1
X_1617_ VGND VDPWR VDPWR VGND _0282_ net91 dig_ctrl_inst.latch_mem_inst.RAM\[41\]\[0\]
+ net119 net53 sky130_fd_sc_hd__and4_1
Xfanout204 VGND VDPWR VDPWR VGND net283 net204 sky130_fd_sc_hd__clkbuf_2
Xfanout226 VGND VDPWR VDPWR VGND net227 net226 sky130_fd_sc_hd__clkbuf_2
Xfanout259 VGND VDPWR VDPWR VGND net259 net260 sky130_fd_sc_hd__buf_1
X_1479_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[0\]\[7\] _0171_ net176
+ _0172_ sky130_fd_sc_hd__o21a_2
Xfanout237 VGND VDPWR VDPWR VGND net237 net244 sky130_fd_sc_hd__buf_1
Xfanout215 VGND VDPWR VDPWR VGND net216 net215 sky130_fd_sc_hd__clkbuf_2
X_1548_ VDPWR VGND VDPWR VGND dig_ctrl_inst.cpu_inst.ip\[4\] _0213_ _0024_ _0197_
+ _0215_ sky130_fd_sc_hd__a22o_1
Xfanout248 VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.instr\[4\] net248 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_49_221 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_32_165 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_305 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_1_3 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_29 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[55\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND net200 dig_ctrl_inst.latch_mem_inst.gclk\[55\] dig_ctrl_inst.latch_mem_inst.RAM\[55\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
X_2451_ VGND VDPWR VDPWR VGND _1032_ _1031_ _1023_ sky130_fd_sc_hd__nand2_1
X_1402_ VGND VDPWR VDPWR VGND _0134_ _1170_ _1156_ sky130_fd_sc_hd__and2b_1
X_2520_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[0\]\[0\] net156 _0046_
+ clknet_leaf_8_clk sky130_fd_sc_hd__dfrtp_4
Xinput4 VGND VDPWR VDPWR VGND net4 ui_in[1] sky130_fd_sc_hd__clkbuf_1
X_1264_ VGND VDPWR VDPWR VGND _1106_ net265 _1092_ _1091_ _1105_ sky130_fd_sc_hd__o31a_2
X_1333_ VGND VDPWR VDPWR VGND _1106_ _1174_ _1052_ _1090_ sky130_fd_sc_hd__nor3_1
X_2382_ VGND VDPWR VDPWR VGND _1003_ _0992_ net342 _0070_ sky130_fd_sc_hd__mux2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[44\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND net213 dig_ctrl_inst.latch_mem_inst.gclk\[44\] dig_ctrl_inst.latch_mem_inst.RAM\[44\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
X_1195_ VDPWR VGND VDPWR VGND net246 _1039_ sky130_fd_sc_hd__inv_2
Xdig_ctrl_inst.latch_mem_inst.genblk1\[2\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[2\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[2\]._gclk clknet_leaf_13_clk sky130_fd_sc_hd__dlclkp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[33\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND net235 dig_ctrl_inst.latch_mem_inst.gclk\[33\] dig_ctrl_inst.latch_mem_inst.RAM\[33\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[25\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[25\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[25\]._gclk clknet_leaf_13_clk sky130_fd_sc_hd__dlclkp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[59\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND net194 dig_ctrl_inst.latch_mem_inst.gclk\[59\] dig_ctrl_inst.latch_mem_inst.RAM\[59\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[10\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND net188 dig_ctrl_inst.latch_mem_inst.gclk\[10\] dig_ctrl_inst.latch_mem_inst.RAM\[10\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
X_1951_ VGND VDPWR VDPWR VGND _0611_ net102 dig_ctrl_inst.latch_mem_inst.RAM\[55\]\[5\]
+ net107 net47 sky130_fd_sc_hd__and4_1
X_1882_ VDPWR VGND VDPWR VGND _0543_ _0126_ dig_ctrl_inst.latch_mem_inst.RAM\[8\]\[4\]
+ dig_ctrl_inst.latch_mem_inst.RAM\[21\]\[4\] _1187_ _0542_ sky130_fd_sc_hd__a221o_1
X_2365_ VDPWR VGND VDPWR VGND _0766_ _0998_ _0946_ _0948_ sky130_fd_sc_hd__o21bai_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[48\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND net203 dig_ctrl_inst.latch_mem_inst.gclk\[48\] dig_ctrl_inst.latch_mem_inst.RAM\[48\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
X_2434_ VDPWR VGND VDPWR VGND dig_ctrl_inst.cpu_inst.cpu_state\[0\] _1015_ _0104_
+ _1021_ _1019_ sky130_fd_sc_hd__a22o_1
X_2503_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.arg1\[0\] net152 _0029_ clknet_leaf_11_clk
+ sky130_fd_sc_hd__dfrtp_1
X_1247_ VDPWR VGND VDPWR VGND net167 net264 _1089_ net166 sky130_fd_sc_hd__a21oi_1
X_1316_ VDPWR VGND VDPWR VGND net252 _1158_ net255 dig_ctrl_inst.cpu_inst.regs\[3\]\[4\]
+ sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[37\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND net225 dig_ctrl_inst.latch_mem_inst.gclk\[37\] dig_ctrl_inst.latch_mem_inst.RAM\[37\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
X_2296_ VGND VDPWR VDPWR VGND _0937_ dig_ctrl_inst.cpu_inst.data\[5\] _0936_ _0813_
+ sky130_fd_sc_hd__a21bo_1
XANTENNA_20 VGND VDPWR VDPWR VGND net327 sky130_fd_sc_hd__diode_2
Xdig_ctrl_inst.latch_mem_inst.genblk1\[38\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[38\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[38\]._gclk sky130_fd_sc_hd__clkbuf_4
X_2607__281 VGND VDPWR VDPWR VGND _2607__281/LO net281 sky130_fd_sc_hd__conb_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[26\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND net243 dig_ctrl_inst.latch_mem_inst.gclk\[26\] dig_ctrl_inst.latch_mem_inst.RAM\[26\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[14\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND net178 dig_ctrl_inst.latch_mem_inst.gclk\[14\] dig_ctrl_inst.latch_mem_inst.RAM\[14\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_0_305 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2081_ VDPWR VGND VDPWR VGND _0739_ _0146_ dig_ctrl_inst.latch_mem_inst.RAM\[40\]\[7\]
+ dig_ctrl_inst.latch_mem_inst.RAM\[43\]\[7\] _0143_ _0738_ sky130_fd_sc_hd__a221o_1
X_2150_ VGND VDPWR VDPWR VGND _0796_ _0794_ _0789_ sky130_fd_sc_hd__nand2_1
X_1934_ VGND VDPWR VDPWR VGND _0594_ net108 dig_ctrl_inst.latch_mem_inst.RAM\[11\]\[5\]
+ net129 net90 sky130_fd_sc_hd__and4_1
XFILLER_0_33_97 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_53 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[8\].gen_latches\[0\].p_latch VGND VDPWR VDPWR
+ VGND net236 dig_ctrl_inst.latch_mem_inst.gclk\[8\] dig_ctrl_inst.latch_mem_inst.RAM\[8\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
X_1865_ VDPWR VGND VDPWR VGND net100 _0526_ dig_ctrl_inst.latch_mem_inst.RAM\[20\]\[4\]
+ net65 sky130_fd_sc_hd__and3_2
X_1796_ VGND VDPWR VDPWR VGND _0456_ _0459_ _0458_ dig_ctrl_inst.latch_mem_inst.RAM\[51\]\[2\]
+ _0153_ _0457_ sky130_fd_sc_hd__a2111o_1
X_2417_ VGND VDPWR VDPWR VGND _0825_ _1013_ _1067_ _0186_ sky130_fd_sc_hd__nor3_1
XPHY_EDGE_ROW_10_Left_88 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2348_ VDPWR VGND VDPWR VGND _0974_ _0987_ _0982_ _0986_ sky130_fd_sc_hd__or3_1
XFILLER_0_66_105 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2279_ VGND VDPWR VDPWR VGND _0915_ _0815_ _0764_ _0921_ sky130_fd_sc_hd__mux2_1
X_1650_ VDPWR VGND VDPWR VGND net87 _0315_ dig_ctrl_inst.latch_mem_inst.RAM\[56\]\[0\]
+ net44 sky130_fd_sc_hd__and3_2
X_1581_ VGND VDPWR VDPWR VGND _0247_ _0246_ _0244_ sky130_fd_sc_hd__nand2_1
X_2202_ VDPWR VGND VDPWR VGND _0847_ _0813_ net160 dig_ctrl_inst.cpu_inst.data\[1\]
+ _0812_ _0846_ sky130_fd_sc_hd__a221o_1
X_2064_ VGND VDPWR VDPWR VGND _0722_ net106 dig_ctrl_inst.latch_mem_inst.RAM\[51\]\[7\]
+ net136 net44 sky130_fd_sc_hd__and4_1
XFILLER_0_44_52 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_2133_ VDPWR VGND VDPWR VGND _0778_ _0779_ sky130_fd_sc_hd__inv_2
X_1917_ VDPWR VGND VDPWR VGND _0270_ _0577_ _0031_ _0576_ sky130_fd_sc_hd__a21oi_1
X_1779_ VDPWR VGND VDPWR VGND _0442_ _0272_ dig_ctrl_inst.latch_mem_inst.RAM\[39\]\[2\]
+ dig_ctrl_inst.latch_mem_inst.RAM\[5\]\[2\] _0142_ _0441_ sky130_fd_sc_hd__a221o_1
X_1848_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[45\]\[3\] _0147_ _0510_
+ dig_ctrl_inst.latch_mem_inst.RAM\[47\]\[3\] _0149_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_290 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_193 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.genblk1\[7\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[7\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[7\]._gclk clknet_leaf_1_clk sky130_fd_sc_hd__dlclkp_1
X_1702_ VGND VDPWR VDPWR VGND _0366_ net77 dig_ctrl_inst.latch_mem_inst.RAM\[63\]\[1\]
+ net110 net44 sky130_fd_sc_hd__and4_1
X_1633_ VDPWR VGND VDPWR VGND _0296_ _0294_ _0298_ _0295_ _0297_ sky130_fd_sc_hd__or4_1
XFILLER_0_5_249 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
X_1564_ VGND VDPWR VDPWR VGND _0227_ _0230_ _0168_ sky130_fd_sc_hd__nor2_1
X_1495_ VGND VDPWR VDPWR VGND _0183_ _0182_ _0180_ dig_ctrl_inst.cpu_inst.data\[1\]
+ dig_ctrl_inst.cpu_inst.data\[0\] sky130_fd_sc_hd__and4b_4
X_2116_ VGND VDPWR VDPWR VGND _1051_ net314 dig_ctrl_inst.cpu_inst.cpu_state\[1\]
+ _0044_ sky130_fd_sc_hd__mux2_1
X_2047_ VGND VDPWR VDPWR VGND _0703_ _0706_ _0705_ dig_ctrl_inst.latch_mem_inst.RAM\[20\]\[6\]
+ _0125_ _0704_ sky130_fd_sc_hd__a2111o_1
Xfanout37 VGND VDPWR VDPWR VGND net42 net37 sky130_fd_sc_hd__clkbuf_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[63\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND net234 dig_ctrl_inst.latch_mem_inst.gclk\[63\] dig_ctrl_inst.latch_mem_inst.RAM\[63\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_44_141 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
Xfanout59 VGND VDPWR VDPWR VGND net61 net59 sky130_fd_sc_hd__clkbuf_2
Xfanout48 VDPWR VGND VDPWR VGND net48 net51 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_13_Left_91 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.genblk1\[32\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[32\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[32\]._gclk clknet_leaf_13_clk sky130_fd_sc_hd__dlclkp_1
Xclkload18 VGND VDPWR VDPWR VGND clknet_leaf_19_clk clkload18/Y sky130_fd_sc_hd__inv_12
X_1280_ VGND VDPWR VDPWR VGND _1121_ _1115_ _1108_ _1044_ _1122_ net265 sky130_fd_sc_hd__a32oi_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[40\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND net187 dig_ctrl_inst.latch_mem_inst.gclk\[40\] dig_ctrl_inst.latch_mem_inst.RAM\[40\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_26_141 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xfanout227 VDPWR VGND VDPWR VGND net227 net285 sky130_fd_sc_hd__buf_2
Xfanout216 VGND VDPWR VDPWR VGND net289 net216 sky130_fd_sc_hd__clkbuf_2
X_2596_ VDPWR VGND VDPWR VGND dig_ctrl_inst.spi_addr\[3\] clknet_leaf_3_clk _0110_
+ sky130_fd_sc_hd__dfxtp_1
Xfanout238 VGND VDPWR VDPWR VGND net241 net238 sky130_fd_sc_hd__clkbuf_2
X_1616_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[8\]\[0\] _1187_ _0281_
+ dig_ctrl_inst.latch_mem_inst.RAM\[40\]\[0\] _0143_ sky130_fd_sc_hd__a22o_1
Xfanout205 VGND VDPWR VDPWR VGND net206 net205 sky130_fd_sc_hd__clkbuf_2
X_1547_ VDPWR VGND VDPWR VGND _1046_ _0209_ _0215_ _0185_ _0214_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_53 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_49_200 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_1478_ VGND VDPWR VDPWR VGND _1063_ _0171_ _0170_ _1038_ dig_ctrl_inst.cpu_inst.regs\[1\]\[7\]
+ _0169_ sky130_fd_sc_hd__a2111o_1
Xfanout249 VGND VDPWR VDPWR VGND net249 net250 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_97 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_233 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_49_277 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_17_174 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_32_177 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_141 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[56\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND net240 dig_ctrl_inst.latch_mem_inst.gclk\[56\] dig_ctrl_inst.latch_mem_inst.RAM\[56\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
X_2381_ VGND VDPWR VDPWR VGND _1066_ _1003_ _0769_ _0189_ sky130_fd_sc_hd__and3b_4
X_2450_ VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_addr\[4\] _1022_ dig_ctrl_inst.spi_addr\[3\]
+ _1027_ _1031_ sky130_fd_sc_hd__a31o_1
X_1401_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[31\] _0133_ _1173_
+ sky130_fd_sc_hd__and2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[0\].gen_latches\[2\].p_latch VGND VDPWR VDPWR
+ VGND net222 dig_ctrl_inst.latch_mem_inst.gclk\[0\] dig_ctrl_inst.latch_mem_inst.RAM\[0\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[44\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND net181 dig_ctrl_inst.latch_mem_inst.gclk\[44\] dig_ctrl_inst.latch_mem_inst.RAM\[44\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
X_1194_ VDPWR VGND VDPWR VGND net251 _1038_ sky130_fd_sc_hd__inv_2
Xinput5 VGND VDPWR VDPWR VGND net5 ui_in[2] sky130_fd_sc_hd__clkbuf_1
X_1263_ VGND VDPWR VDPWR VGND _1105_ _1098_ _1082_ _1104_ _1055_ _1070_ sky130_fd_sc_hd__a32o_1
X_1332_ VDPWR VGND VDPWR VGND net126 dig_ctrl_inst.latch_mem_inst.data_we\[0\] net133
+ _1173_ sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[33\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND net201 dig_ctrl_inst.latch_mem_inst.gclk\[33\] dig_ctrl_inst.latch_mem_inst.RAM\[33\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_72_3 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2579_ VGND VDPWR VDPWR VGND net30 net172 _0093_ clknet_leaf_5_clk sky130_fd_sc_hd__dfrtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[22\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND net216 dig_ctrl_inst.latch_mem_inst.gclk\[22\] dig_ctrl_inst.latch_mem_inst.RAM\[22\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_20_158 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_29_Left_107 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[11\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND net231 dig_ctrl_inst.latch_mem_inst.gclk\[11\] dig_ctrl_inst.latch_mem_inst.RAM\[11\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_38_Left_116 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_7_108 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1950_ VDPWR VGND VDPWR VGND net111 _0610_ dig_ctrl_inst.latch_mem_inst.RAM\[18\]\[5\]
+ net59 sky130_fd_sc_hd__and3_2
X_1881_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[7\]\[4\] _1184_ _0542_
+ dig_ctrl_inst.latch_mem_inst.RAM\[59\]\[4\] _0159_ sky130_fd_sc_hd__a22o_1
X_2502_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.arg0\[1\] net154 _0028_ clknet_leaf_11_clk
+ sky130_fd_sc_hd__dfrtp_1
X_2364_ VGND VDPWR VDPWR VGND _0991_ _0997_ net340 _0058_ sky130_fd_sc_hd__mux2_1
X_2433_ VGND VDPWR VDPWR VGND _1020_ _1021_ _1015_ sky130_fd_sc_hd__nor2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[4\].gen_latches\[3\].p_latch VGND VDPWR VDPWR
+ VGND net217 dig_ctrl_inst.latch_mem_inst.gclk\[4\] dig_ctrl_inst.latch_mem_inst.RAM\[4\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_47_Left_125 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1315_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.ip\[4\] _1073_ _1071_ _1053_
+ _1157_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_56_Left_134 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1246_ VDPWR VGND VDPWR VGND net165 _1088_ sky130_fd_sc_hd__inv_2
X_2295_ VGND VDPWR VDPWR VGND _0806_ _0936_ _0810_ _1147_ _0930_ sky130_fd_sc_hd__o22a_1
XANTENNA_10 VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[24\] sky130_fd_sc_hd__diode_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[37\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND net190 dig_ctrl_inst.latch_mem_inst.gclk\[37\] dig_ctrl_inst.latch_mem_inst.RAM\[37\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
XANTENNA_21 VGND VDPWR VDPWR VGND _0461_ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_65_Left_143 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_74_Left_152 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[26\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND net207 dig_ctrl_inst.latch_mem_inst.gclk\[26\] dig_ctrl_inst.latch_mem_inst.RAM\[26\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[15\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND net223 dig_ctrl_inst.latch_mem_inst.gclk\[15\] dig_ctrl_inst.latch_mem_inst.RAM\[15\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_68_29 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_48_309 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2080_ VGND VDPWR VDPWR VGND _0738_ net60 dig_ctrl_inst.latch_mem_inst.RAM\[46\]\[7\]
+ _0148_ dig_ctrl_inst.latch_mem_inst.RAM\[24\]\[7\] net85 sky130_fd_sc_hd__a32o_1
X_1933_ VDPWR VGND VDPWR VGND net81 _0593_ dig_ctrl_inst.latch_mem_inst.RAM\[26\]\[5\]
+ net63 sky130_fd_sc_hd__and3_2
X_1864_ VDPWR VGND VDPWR VGND net128 _0525_ dig_ctrl_inst.latch_mem_inst.RAM\[4\]\[4\]
+ net100 sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[8\].gen_latches\[4\].p_latch VGND VDPWR VDPWR
+ VGND net208 dig_ctrl_inst.latch_mem_inst.gclk\[8\] dig_ctrl_inst.latch_mem_inst.RAM\[8\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
X_1795_ VDPWR VGND VDPWR VGND net73 _0458_ dig_ctrl_inst.latch_mem_inst.RAM\[60\]\[2\]
+ net45 sky130_fd_sc_hd__and3_2
XFILLER_0_31_209 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
X_2416_ VGND VDPWR VDPWR VGND _1012_ dig_ctrl_inst.cpu_inst.port_o\[7\] net32 _0095_
+ sky130_fd_sc_hd__mux2_1
X_2347_ VGND VDPWR VDPWR VGND _0884_ _0986_ _0984_ _1114_ net162 _0985_ sky130_fd_sc_hd__o221a_1
X_2278_ VGND VDPWR VDPWR VGND _0919_ _0917_ _0810_ _0234_ _0920_ sky130_fd_sc_hd__o211a_1
X_1229_ VGND VDPWR VDPWR VGND net177 _1062_ net176 _1060_ _1071_ _1057_ sky130_fd_sc_hd__o32ai_4
Xdig_ctrl_inst.latch_mem_inst.genblk1\[37\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[37\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[37\]._gclk clknet_leaf_1_clk sky130_fd_sc_hd__dlclkp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[19\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND net216 dig_ctrl_inst.latch_mem_inst.gclk\[19\] dig_ctrl_inst.latch_mem_inst.RAM\[19\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_53_323 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1580_ VGND VDPWR VDPWR VGND _1129_ _0246_ net160 sky130_fd_sc_hd__or2_1
XFILLER_0_0_103 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_0_169 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_2201_ VGND VDPWR VDPWR VGND _0810_ _0846_ _0262_ sky130_fd_sc_hd__nor2_1
X_2132_ VGND VDPWR VDPWR VGND _0778_ net140 net159 sky130_fd_sc_hd__nand2_1
X_2063_ VDPWR VGND VDPWR VGND net81 _0721_ dig_ctrl_inst.latch_mem_inst.RAM\[58\]\[7\]
+ net44 sky130_fd_sc_hd__and3_2
X_1847_ VGND VDPWR VDPWR VGND _0479_ _0509_ _0489_ dig_ctrl_inst.latch_mem_inst.RAM\[23\]\[3\]
+ _0128_ _0486_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_8_236 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_1916_ VGND VDPWR VDPWR VGND _0270_ _0577_ net248 sky130_fd_sc_hd__nor2_1
X_1778_ VDPWR VGND VDPWR VGND net74 _0441_ dig_ctrl_inst.latch_mem_inst.RAM\[44\]\[2\]
+ net55 sky130_fd_sc_hd__and3_2
XFILLER_0_69_50 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
X_1701_ VGND VDPWR VDPWR VGND _0364_ _0357_ _0365_ _0345_ _0350_ sky130_fd_sc_hd__nor4_1
X_1632_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[18\]\[0\] _0123_ _0297_
+ dig_ctrl_inst.latch_mem_inst.RAM\[55\]\[0\] _0155_ sky130_fd_sc_hd__a22o_1
X_1563_ VDPWR VGND VDPWR VGND _0228_ _0229_ sky130_fd_sc_hd__inv_2
X_1494_ VDPWR VGND VDPWR VGND _0181_ _0182_ sky130_fd_sc_hd__inv_2
X_2115_ VGND VDPWR VDPWR VGND _1051_ net313 dig_ctrl_inst.cpu_inst.cpu_state\[0\]
+ _0043_ sky130_fd_sc_hd__mux2_1
X_2046_ VDPWR VGND VDPWR VGND _1177_ _0705_ dig_ctrl_inst.latch_mem_inst.RAM\[18\]\[6\]
+ net66 sky130_fd_sc_hd__and3_2
Xfanout49 VGND VDPWR VDPWR VGND net49 net51 sky130_fd_sc_hd__buf_1
Xfanout38 VDPWR VGND VDPWR VGND net42 net38 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_44_153 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
Xdig_ctrl_inst.latch_mem_inst.gen_words\[63\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND net202 dig_ctrl_inst.latch_mem_inst.gclk\[63\] dig_ctrl_inst.latch_mem_inst.RAM\[63\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[52\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND net218 dig_ctrl_inst.latch_mem_inst.gclk\[52\] dig_ctrl_inst.latch_mem_inst.RAM\[52\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_35_120 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_50_189 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
Xdig_ctrl_inst.latch_mem_inst.gen_words\[41\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND net228 dig_ctrl_inst.latch_mem_inst.gclk\[41\] dig_ctrl_inst.latch_mem_inst.RAM\[41\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_18_109 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1477_ VGND VDPWR VDPWR VGND net255 net251 _0170_ dig_ctrl_inst.cpu_inst.regs\[2\]\[7\]
+ sky130_fd_sc_hd__and3b_1
Xfanout217 VGND VDPWR VDPWR VGND net218 net217 sky130_fd_sc_hd__clkbuf_2
X_2595_ VDPWR VGND VDPWR VGND dig_ctrl_inst.spi_addr\[2\] clknet_leaf_3_clk _0109_
+ sky130_fd_sc_hd__dfxtp_1
X_1615_ VGND VDPWR VDPWR VGND _0280_ net62 dig_ctrl_inst.latch_mem_inst.RAM\[38\]\[0\]
+ _0141_ dig_ctrl_inst.latch_mem_inst.RAM\[28\]\[0\] net72 sky130_fd_sc_hd__a32o_1
Xfanout228 VGND VDPWR VDPWR VGND net229 net228 sky130_fd_sc_hd__clkbuf_2
X_1546_ VGND VDPWR VDPWR VGND _0191_ net158 dig_ctrl_inst.cpu_inst.data\[4\] _0214_
+ sky130_fd_sc_hd__mux2_1
Xfanout206 VGND VDPWR VDPWR VGND net283 net206 sky130_fd_sc_hd__clkbuf_2
Xfanout239 VGND VDPWR VDPWR VGND net239 net241 sky130_fd_sc_hd__buf_1
X_2029_ VGND VDPWR VDPWR VGND _0688_ net120 dig_ctrl_inst.latch_mem_inst.RAM\[17\]\[6\]
+ net136 net67 sky130_fd_sc_hd__and4_1
XFILLER_0_17_164 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_32_189 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
Xdig_ctrl_inst.latch_mem_inst.gen_words\[56\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND net204 dig_ctrl_inst.latch_mem_inst.gclk\[56\] dig_ctrl_inst.latch_mem_inst.RAM\[56\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[41\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[41\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[41\]._gclk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_63_281 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[45\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND net225 dig_ctrl_inst.latch_mem_inst.gclk\[45\] dig_ctrl_inst.latch_mem_inst.RAM\[45\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_23_101 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_23_123 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2380_ VGND VDPWR VDPWR VGND _1002_ _1001_ net333 _0069_ sky130_fd_sc_hd__mux2_1
X_1331_ VGND VDPWR VDPWR VGND _1173_ net167 dig_ctrl_inst.mode_sync dig_ctrl_inst.spi_receiver_inst.stb_o
+ sky130_fd_sc_hd__a21o_2
X_1400_ VDPWR VGND VDPWR VGND net76 _0133_ net105 net62 sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[34\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND net241 dig_ctrl_inst.latch_mem_inst.gclk\[34\] dig_ctrl_inst.latch_mem_inst.RAM\[34\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
Xinput6 VGND VDPWR VDPWR VGND net6 ui_in[3] sky130_fd_sc_hd__clkbuf_1
X_1193_ VDPWR VGND VDPWR VGND dig_ctrl_inst.cpu_inst.cpu_state\[1\] _1037_ sky130_fd_sc_hd__inv_2
X_1262_ VGND VDPWR VDPWR VGND net177 _1100_ _1101_ _1102_ _1103_ _1104_ sky130_fd_sc_hd__o41a_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[0\].gen_latches\[6\].p_latch VGND VDPWR VDPWR
+ VGND net284 dig_ctrl_inst.latch_mem_inst.gclk\[0\] dig_ctrl_inst.latch_mem_inst.RAM\[0\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_46_248 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2578_ VGND VDPWR VDPWR VGND net29 net172 _0092_ clknet_leaf_6_clk sky130_fd_sc_hd__dfrtp_1
X_1529_ VGND VDPWR VDPWR VGND _0200_ dig_ctrl_inst.cpu_inst.ip\[1\] dig_ctrl_inst.cpu_inst.ip\[0\]
+ sky130_fd_sc_hd__nand2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[22\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND net185 dig_ctrl_inst.latch_mem_inst.gclk\[22\] dig_ctrl_inst.latch_mem_inst.RAM\[22\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_45_281 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_14_Right_14 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[11\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND net201 dig_ctrl_inst.latch_mem_inst.gclk\[11\] dig_ctrl_inst.latch_mem_inst.RAM\[11\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_23_Right_23 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.genblk1\[44\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[44\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[44\]._gclk clknet_leaf_16_clk sky130_fd_sc_hd__dlclkp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[49\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND net215 dig_ctrl_inst.latch_mem_inst.gclk\[49\] dig_ctrl_inst.latch_mem_inst.RAM\[49\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
X_1880_ VGND VDPWR VDPWR VGND _0541_ net88 dig_ctrl_inst.latch_mem_inst.RAM\[43\]\[4\]
+ net104 net50 sky130_fd_sc_hd__and4_1
XFILLER_0_28_204 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_32_Right_32 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_3_337 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2501_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.arg0\[0\] net153 _0027_ clknet_leaf_11_clk
+ sky130_fd_sc_hd__dfrtp_1
X_1314_ VDPWR VGND VDPWR VGND _1156_ _1155_ _1142_ _1154_ dig_ctrl_inst.spi_addr\[5\]
+ _1041_ sky130_fd_sc_hd__o32a_1
X_2363_ VDPWR VGND VDPWR VGND _0766_ _0997_ _0923_ _0926_ sky130_fd_sc_hd__o21bai_1
XPHY_EDGE_ROW_41_Right_41 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[38\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND net231 dig_ctrl_inst.latch_mem_inst.gclk\[38\] dig_ctrl_inst.latch_mem_inst.RAM\[38\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
X_2294_ VGND VDPWR VDPWR VGND _0913_ _0935_ net159 sky130_fd_sc_hd__xnor2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[4\].gen_latches\[7\].p_latch VGND VDPWR VDPWR
+ VGND net180 dig_ctrl_inst.latch_mem_inst.gclk\[4\] dig_ctrl_inst.latch_mem_inst.RAM\[4\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
X_2432_ VGND VDPWR VDPWR VGND _0189_ net248 _1020_ dig_ctrl_inst.cpu_inst.instr\[5\]
+ _1059_ sky130_fd_sc_hd__and4b_1
XPHY_EDGE_ROW_50_Right_50 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1245_ VGND VDPWR VDPWR VGND net177 _1083_ _1084_ _1085_ _1086_ _1087_ sky130_fd_sc_hd__o41a_1
XFILLER_0_63_52 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XANTENNA_11 VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[24\] sky130_fd_sc_hd__diode_2
XANTENNA_22 VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[44\] sky130_fd_sc_hd__diode_2
XFILLER_0_6_120 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_6_197 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_33_240 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[15\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND net186 dig_ctrl_inst.latch_mem_inst.gclk\[15\] dig_ctrl_inst.latch_mem_inst.RAM\[15\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
X_1863_ VDPWR VGND VDPWR VGND net73 _0524_ dig_ctrl_inst.latch_mem_inst.RAM\[28\]\[4\]
+ net64 sky130_fd_sc_hd__and3_2
X_1932_ VDPWR VGND VDPWR VGND net81 _0592_ dig_ctrl_inst.latch_mem_inst.RAM\[42\]\[5\]
+ net55 sky130_fd_sc_hd__and3_2
X_2415_ VGND VDPWR VDPWR VGND _1012_ dig_ctrl_inst.cpu_inst.port_o\[6\] net31 _0094_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_41 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1794_ VDPWR VGND VDPWR VGND net130 _0457_ dig_ctrl_inst.latch_mem_inst.RAM\[8\]\[2\]
+ net86 sky130_fd_sc_hd__and3_2
XFILLER_0_58_85 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_28_3 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_2346_ VGND VDPWR VDPWR VGND _0985_ _0983_ _0909_ _0794_ _0887_ sky130_fd_sc_hd__a211o_1
X_2277_ VGND VDPWR VDPWR VGND _0919_ _0918_ _1162_ _0807_ net159 _0812_ sky130_fd_sc_hd__a221oi_1
X_1228_ VGND VDPWR VDPWR VGND _1060_ _1057_ net176 _1062_ net177 _1070_ sky130_fd_sc_hd__o32a_2
Xdig_ctrl_inst.latch_mem_inst.genblk1\[34\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[34\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[34\]._gclk sky130_fd_sc_hd__clkbuf_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[19\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND net178 dig_ctrl_inst.latch_mem_inst.gclk\[19\] dig_ctrl_inst.latch_mem_inst.RAM\[19\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
X_2062_ VDPWR VGND VDPWR VGND net84 _0720_ dig_ctrl_inst.latch_mem_inst.RAM\[56\]\[7\]
+ net37 sky130_fd_sc_hd__and3_2
X_2131_ VGND VDPWR VDPWR VGND _0172_ _0168_ _0777_ _1147_ _1162_ sky130_fd_sc_hd__nor4_1
X_2200_ VGND VDPWR VDPWR VGND _0844_ _1098_ _0806_ _0845_ net165 sky130_fd_sc_hd__a2bb2o_1
X_1846_ VGND VDPWR VDPWR VGND _0485_ _0508_ _0507_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_248 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1915_ VGND VDPWR VDPWR VGND _0576_ _0575_ _0574_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_14_clk VGND VDPWR VDPWR VGND clknet_leaf_14_clk clknet_1_0__leaf_clk
+ sky130_fd_sc_hd__clkbuf_8
X_1777_ VGND VDPWR VDPWR VGND _0437_ _0440_ _0439_ dig_ctrl_inst.latch_mem_inst.RAM\[9\]\[2\]
+ _1188_ _0438_ sky130_fd_sc_hd__a2111o_1
XPHY_EDGE_ROW_4_Right_4 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_39_107 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2329_ VGND VDPWR VDPWR VGND _0227_ _0969_ _0947_ sky130_fd_sc_hd__or2_1
XFILLER_0_53_143 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_1631_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[16\]\[0\] _0121_ _0296_
+ dig_ctrl_inst.latch_mem_inst.RAM\[5\]\[0\] _0272_ sky130_fd_sc_hd__a22o_1
X_1700_ VDPWR VGND VDPWR VGND _0358_ _0364_ _0359_ _0363_ sky130_fd_sc_hd__or3_1
Xclkbuf_leaf_3_clk VGND VDPWR VDPWR VGND clknet_leaf_3_clk clknet_1_1__leaf_clk sky130_fd_sc_hd__clkbuf_8
X_1562_ VDPWR VGND VDPWR VGND _0228_ _0227_ _0168_ sky130_fd_sc_hd__and2_1
X_1493_ VDPWR VGND VDPWR VGND dig_ctrl_inst.cpu_inst.data\[7\] dig_ctrl_inst.cpu_inst.data\[5\]
+ _0181_ dig_ctrl_inst.cpu_inst.data\[4\] dig_ctrl_inst.cpu_inst.data\[6\] sky130_fd_sc_hd__or4_1
X_2045_ VDPWR VGND VDPWR VGND net82 _0704_ dig_ctrl_inst.latch_mem_inst.RAM\[26\]\[6\]
+ net66 sky130_fd_sc_hd__and3_2
XFILLER_0_55_97 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2114_ VGND VDPWR VDPWR VGND _0762_ _0761_ net329 _0042_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_41 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
Xfanout39 VDPWR VGND VDPWR VGND net39 net42 sky130_fd_sc_hd__buf_2
X_1829_ VDPWR VGND VDPWR VGND net129 _0491_ dig_ctrl_inst.latch_mem_inst.RAM\[4\]\[3\]
+ net98 sky130_fd_sc_hd__and3_2
Xmax_cap161 VGND VDPWR VDPWR VGND net162 net161 sky130_fd_sc_hd__clkbuf_2
Xdig_ctrl_inst.latch_mem_inst.genblk1\[49\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[49\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[49\]._gclk clknet_leaf_19_clk sky130_fd_sc_hd__dlclkp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[52\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND net183 dig_ctrl_inst.latch_mem_inst.gclk\[52\] dig_ctrl_inst.latch_mem_inst.RAM\[52\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_35_132 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
Xdig_ctrl_inst.latch_mem_inst.gen_words\[41\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND net195 dig_ctrl_inst.latch_mem_inst.gclk\[41\] dig_ctrl_inst.latch_mem_inst.RAM\[41\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[51\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[51\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[51\]._gclk clknet_leaf_1_clk sky130_fd_sc_hd__dlclkp_1
XFILLER_0_41_22 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[30\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND net217 dig_ctrl_inst.latch_mem_inst.gclk\[30\] dig_ctrl_inst.latch_mem_inst.RAM\[30\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
X_2594_ VDPWR VGND VDPWR VGND dig_ctrl_inst.spi_addr\[1\] clknet_leaf_3_clk _0108_
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_113 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1614_ VDPWR VGND VDPWR VGND _0277_ _0279_ _0271_ sky130_fd_sc_hd__or2_2
Xfanout218 VGND VDPWR VDPWR VGND net289 net218 sky130_fd_sc_hd__clkbuf_2
X_1476_ VDPWR VGND VDPWR VGND net251 _0169_ net255 dig_ctrl_inst.cpu_inst.regs\[3\]\[7\]
+ sky130_fd_sc_hd__and3_2
Xfanout207 VGND VDPWR VDPWR VGND net208 net207 sky130_fd_sc_hd__clkbuf_2
Xfanout229 VGND VDPWR VDPWR VGND net230 net229 sky130_fd_sc_hd__clkbuf_2
X_1545_ VGND VDPWR VDPWR VGND _0213_ _0212_ _0197_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_33 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2028_ VGND VDPWR VDPWR VGND _0687_ net78 dig_ctrl_inst.latch_mem_inst.RAM\[61\]\[6\]
+ net120 net45 sky130_fd_sc_hd__and4_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[27\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[27\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[27\]._gclk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_47 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_11_308 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
Xdig_ctrl_inst.latch_mem_inst.gen_words\[1\].gen_latches\[1\].p_latch VGND VDPWR VDPWR
+ VGND net233 dig_ctrl_inst.latch_mem_inst.gclk\[1\] dig_ctrl_inst.latch_mem_inst.RAM\[1\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
X_1330_ VDPWR VGND VDPWR VGND net128 _1172_ sky130_fd_sc_hd__inv_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[45\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND net194 dig_ctrl_inst.latch_mem_inst.gclk\[45\] dig_ctrl_inst.latch_mem_inst.RAM\[45\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
X_1261_ VDPWR VGND VDPWR VGND net261 _1103_ net257 dig_ctrl_inst.cpu_inst.regs\[0\]\[1\]
+ sky130_fd_sc_hd__or3_1
X_1192_ VDPWR VGND VDPWR VGND dig_ctrl_inst.cpu_inst.cpu_state\[0\] _1036_ sky130_fd_sc_hd__inv_2
Xinput7 VGND VDPWR VDPWR VGND net7 ui_in[4] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_99 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[34\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND net204 dig_ctrl_inst.latch_mem_inst.gclk\[34\] dig_ctrl_inst.latch_mem_inst.RAM\[34\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
X_2577_ VGND VDPWR VDPWR VGND net28 net172 _0091_ clknet_leaf_6_clk sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_3 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
Xdig_ctrl_inst.latch_mem_inst.gen_words\[23\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND net226 dig_ctrl_inst.latch_mem_inst.gclk\[23\] dig_ctrl_inst.latch_mem_inst.RAM\[23\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_77_51 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1459_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[61\] _0161_ net147
+ sky130_fd_sc_hd__and2_1
X_1528_ VGND VDPWR VDPWR VGND _0197_ _0199_ dig_ctrl_inst.cpu_inst.ip\[0\] _0020_
+ sky130_fd_sc_hd__mux2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[12\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND net243 dig_ctrl_inst.latch_mem_inst.gclk\[12\] dig_ctrl_inst.latch_mem_inst.RAM\[12\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[5\].gen_latches\[2\].p_latch VGND VDPWR VDPWR
+ VGND net224 dig_ctrl_inst.latch_mem_inst.gclk\[5\] dig_ctrl_inst.latch_mem_inst.RAM\[5\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[49\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND net182 dig_ctrl_inst.latch_mem_inst.gclk\[49\] dig_ctrl_inst.latch_mem_inst.RAM\[49\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_22_24 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_28_216 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_36_260 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2500_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.skip net152 _0026_ clknet_leaf_14_clk
+ sky130_fd_sc_hd__dfrtp_2
X_2431_ VGND VDPWR VDPWR VGND _1019_ _1016_ _1017_ _0576_ _1018_ sky130_fd_sc_hd__a211o_1
X_1313_ VGND VDPWR VDPWR VGND _1070_ net265 _1055_ _1147_ _1155_ sky130_fd_sc_hd__a31o_1
X_1244_ VDPWR VGND VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[0\]\[0\] _1086_ net262
+ net258 sky130_fd_sc_hd__or3_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[38\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND net200 dig_ctrl_inst.latch_mem_inst.gclk\[38\] dig_ctrl_inst.latch_mem_inst.RAM\[38\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
X_2293_ VGND VDPWR VDPWR VGND _0934_ _0913_ _1153_ sky130_fd_sc_hd__nand2_1
X_2362_ VGND VDPWR VDPWR VGND _0991_ _0996_ net348 _0057_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_20 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_23 VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[52\] sky130_fd_sc_hd__diode_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[27\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND net212 dig_ctrl_inst.latch_mem_inst.gclk\[27\] dig_ctrl_inst.latch_mem_inst.RAM\[27\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
XANTENNA_12 VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[24\] sky130_fd_sc_hd__diode_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[16\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND net235 dig_ctrl_inst.latch_mem_inst.gclk\[16\] dig_ctrl_inst.latch_mem_inst.RAM\[16\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
X_2614__277 VGND VDPWR VDPWR VGND net277 _2614__277/HI sky130_fd_sc_hd__conb_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[9\].gen_latches\[3\].p_latch VGND VDPWR VDPWR
+ VGND net211 dig_ctrl_inst.latch_mem_inst.gclk\[9\] dig_ctrl_inst.latch_mem_inst.RAM\[9\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[7\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[7\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[7\]._gclk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_33_23 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_68_193 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xinput10 VGND VDPWR VDPWR VGND net10 ui_in[7] sky130_fd_sc_hd__clkbuf_1
X_1931_ VDPWR VGND VDPWR VGND net86 _0591_ dig_ctrl_inst.latch_mem_inst.RAM\[40\]\[5\]
+ net53 sky130_fd_sc_hd__and3_2
X_1793_ VGND VDPWR VDPWR VGND _0456_ net79 dig_ctrl_inst.latch_mem_inst.RAM\[29\]\[2\]
+ net120 net66 sky130_fd_sc_hd__and4_1
X_1862_ VGND VDPWR VDPWR VGND _0270_ _0522_ net249 _0030_ sky130_fd_sc_hd__mux2_1
X_2414_ VGND VDPWR VDPWR VGND _1012_ dig_ctrl_inst.cpu_inst.port_o\[5\] net358 _0093_
+ sky130_fd_sc_hd__mux2_1
X_1227_ VDPWR VGND VDPWR VGND _1069_ net260 _1035_ sky130_fd_sc_hd__and2_1
X_2345_ VGND VDPWR VDPWR VGND _0942_ _0984_ _0857_ sky130_fd_sc_hd__nor2_1
X_2276_ VGND VDPWR VDPWR VGND _0817_ _1162_ _0806_ _0918_ _0236_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_47_333 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.genblk1\[56\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[56\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[56\]._gclk clknet_leaf_16_clk sky130_fd_sc_hd__dlclkp_1
X_2130_ VDPWR VGND VDPWR VGND _0775_ _0776_ _1098_ sky130_fd_sc_hd__or2_2
X_2061_ VDPWR VGND VDPWR VGND net125 _0719_ dig_ctrl_inst.latch_mem_inst.RAM\[6\]\[7\]
+ net93 sky130_fd_sc_hd__and3_2
X_1914_ VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[0\]\[4\] _0575_ _0279_
+ sky130_fd_sc_hd__or2_1
X_1845_ VGND VDPWR VDPWR VGND _0507_ net95 dig_ctrl_inst.latch_mem_inst.RAM\[33\]\[3\]
+ _0136_ dig_ctrl_inst.latch_mem_inst.RAM\[6\]\[3\] net129 sky130_fd_sc_hd__a32o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[60\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND net211 dig_ctrl_inst.latch_mem_inst.gclk\[60\] dig_ctrl_inst.latch_mem_inst.RAM\[60\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
X_1776_ VDPWR VGND VDPWR VGND net126 _0439_ dig_ctrl_inst.latch_mem_inst.RAM\[4\]\[2\]
+ net97 sky130_fd_sc_hd__and3_2
X_2328_ VGND VDPWR VDPWR VGND _0968_ _0947_ _0227_ sky130_fd_sc_hd__nand2_1
X_2259_ VDPWR VGND VDPWR VGND _0900_ _0888_ _0902_ _0891_ _0901_ sky130_fd_sc_hd__or4_1
XFILLER_0_38_141 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_53_188 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1630_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[46\]\[0\] _0148_ _0295_
+ dig_ctrl_inst.latch_mem_inst.RAM\[59\]\[0\] _0159_ sky130_fd_sc_hd__a22o_1
X_1561_ VDPWR VGND VDPWR VGND _0227_ net177 _0226_ dig_ctrl_inst.cpu_inst.regs\[0\]\[6\]
+ sky130_fd_sc_hd__mux2_4
X_1492_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.data\[2\] _0180_ dig_ctrl_inst.cpu_inst.data\[3\]
+ sky130_fd_sc_hd__nor2_1
X_2044_ VDPWR VGND VDPWR VGND net99 _0703_ dig_ctrl_inst.latch_mem_inst.RAM\[52\]\[6\]
+ net45 sky130_fd_sc_hd__and3_2
X_2113_ VGND VDPWR VDPWR VGND _0762_ _0709_ net336 _0041_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_185 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1828_ VDPWR VGND VDPWR VGND net94 _0490_ dig_ctrl_inst.latch_mem_inst.RAM\[22\]\[3\]
+ net64 sky130_fd_sc_hd__and3_2
Xmax_cap140 VGND VDPWR VDPWR VGND _0777_ net140 sky130_fd_sc_hd__clkbuf_2
X_1759_ VGND VDPWR VDPWR VGND _0422_ net88 dig_ctrl_inst.latch_mem_inst.RAM\[57\]\[2\]
+ net116 net38 sky130_fd_sc_hd__and4_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[53\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND net227 dig_ctrl_inst.latch_mem_inst.gclk\[53\] dig_ctrl_inst.latch_mem_inst.RAM\[53\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[42\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND net244 dig_ctrl_inst.latch_mem_inst.gclk\[42\] dig_ctrl_inst.latch_mem_inst.RAM\[42\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_25_57 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_25_46 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_26_133 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_41_169 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
Xdig_ctrl_inst.latch_mem_inst.gen_words\[30\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND net184 dig_ctrl_inst.latch_mem_inst.gclk\[30\] dig_ctrl_inst.latch_mem_inst.RAM\[30\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
X_2593_ VDPWR VGND VDPWR VGND dig_ctrl_inst.spi_addr\[0\] clknet_leaf_3_clk _0107_
+ sky130_fd_sc_hd__dfxtp_1
X_1613_ VGND VDPWR VDPWR VGND _0277_ _0278_ _0271_ sky130_fd_sc_hd__nor2_1
X_1544_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.ip\[4\] _0185_ dig_ctrl_inst.cpu_inst.ip\[3\]
+ _0204_ _0212_ sky130_fd_sc_hd__a31o_1
X_1475_ VDPWR VGND VDPWR VGND net266 dig_ctrl_inst.spi_data_o\[6\] dig_ctrl_inst.data_out\[6\]
+ _0168_ _0164_ sky130_fd_sc_hd__a22o_1
X_2601__268 VGND VDPWR VDPWR VGND net268 _2601__268/HI sky130_fd_sc_hd__conb_1
Xfanout208 VDPWR VGND VDPWR VGND net209 net208 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout219 VGND VDPWR VDPWR VGND net220 net219 sky130_fd_sc_hd__clkbuf_2
X_2027_ VDPWR VGND VDPWR VGND net99 _0686_ dig_ctrl_inst.latch_mem_inst.RAM\[36\]\[6\]
+ net55 sky130_fd_sc_hd__and3_2
XFILLER_0_32_103 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_17_Left_95 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[57\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND net216 dig_ctrl_inst.latch_mem_inst.gclk\[57\] dig_ctrl_inst.latch_mem_inst.RAM\[57\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[46\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND net234 dig_ctrl_inst.latch_mem_inst.gclk\[46\] dig_ctrl_inst.latch_mem_inst.RAM\[46\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
Xinput8 VGND VDPWR VDPWR VGND net8 ui_in[5] sky130_fd_sc_hd__clkbuf_1
X_1191_ VDPWR VGND VDPWR VGND net262 _1035_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_23 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1260_ VGND VDPWR VDPWR VGND _1102_ net261 dig_ctrl_inst.cpu_inst.regs\[2\]\[1\]
+ sky130_fd_sc_hd__and2b_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[1\].gen_latches\[5\].p_latch VGND VDPWR VDPWR
+ VGND net197 dig_ctrl_inst.latch_mem_inst.gclk\[1\] dig_ctrl_inst.latch_mem_inst.RAM\[1\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_36_78 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
X_2576_ VGND VDPWR VDPWR VGND net27 net173 _0090_ clknet_leaf_6_clk sky130_fd_sc_hd__dfrtp_1
X_1527_ VGND VDPWR VDPWR VGND _0185_ _0198_ _1040_ _0199_ sky130_fd_sc_hd__mux2_1
X_1458_ VDPWR VGND VDPWR VGND net78 _0161_ net121 net46 sky130_fd_sc_hd__and3_2
X_1389_ VDPWR VGND VDPWR VGND net85 dig_ctrl_inst.latch_mem_inst.data_we\[24\] net143
+ net59 sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[23\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND net186 dig_ctrl_inst.latch_mem_inst.gclk\[23\] dig_ctrl_inst.latch_mem_inst.RAM\[23\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_9_152 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_20_117 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
Xdig_ctrl_inst.latch_mem_inst.gen_words\[12\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND net203 dig_ctrl_inst.latch_mem_inst.gclk\[12\] dig_ctrl_inst.latch_mem_inst.RAM\[12\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[39\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND net243 dig_ctrl_inst.latch_mem_inst.gclk\[39\] dig_ctrl_inst.latch_mem_inst.RAM\[39\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[5\].gen_latches\[6\].p_latch VGND VDPWR VDPWR
+ VGND net190 dig_ctrl_inst.latch_mem_inst.gclk\[5\] dig_ctrl_inst.latch_mem_inst.RAM\[5\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
X_2430_ VGND VDPWR VDPWR VGND _0575_ _0522_ _1018_ _0648_ _0574_ sky130_fd_sc_hd__and4b_1
X_2361_ VDPWR VGND VDPWR VGND _0766_ _0996_ _0902_ _0903_ sky130_fd_sc_hd__o21bai_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[63\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[63\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[63\]._gclk clknet_leaf_15_clk sky130_fd_sc_hd__dlclkp_1
X_1312_ VDPWR VGND VDPWR VGND _1154_ net159 net167 sky130_fd_sc_hd__and2_1
X_1243_ VGND VDPWR VDPWR VGND _1085_ net258 dig_ctrl_inst.cpu_inst.regs\[1\]\[0\]
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_63_32 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_2292_ VGND VDPWR VDPWR VGND _0933_ _0234_ _0931_ _0907_ sky130_fd_sc_hd__nand3_1
XFILLER_0_59_331 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_25_Left_103 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XANTENNA_13 VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[36\] sky130_fd_sc_hd__diode_2
XANTENNA_24 VGND VDPWR VDPWR VGND net28 sky130_fd_sc_hd__diode_2
XFILLER_0_70_3 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_34_209 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2559_ VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_data_o\[3\] net175 _0083_ clknet_leaf_9_clk
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_34_Left_112 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[27\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND net180 dig_ctrl_inst.latch_mem_inst.gclk\[27\] dig_ctrl_inst.latch_mem_inst.RAM\[27\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_43_Left_121 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[16\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND net195 dig_ctrl_inst.latch_mem_inst.gclk\[16\] dig_ctrl_inst.latch_mem_inst.RAM\[16\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_52_Left_130 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_0_309 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_1930_ VGND VDPWR VDPWR VGND _0590_ net79 dig_ctrl_inst.latch_mem_inst.RAM\[30\]\[5\]
+ net115 net67 sky130_fd_sc_hd__and4_1
Xinput11 VGND VDPWR VDPWR VGND net11 uio_in[0] sky130_fd_sc_hd__clkbuf_1
X_1792_ VGND VDPWR VDPWR VGND _0452_ _0455_ _0454_ dig_ctrl_inst.latch_mem_inst.RAM\[30\]\[2\]
+ _0132_ _0453_ sky130_fd_sc_hd__a2111o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[9\].gen_latches\[7\].p_latch VGND VDPWR VDPWR
+ VGND net185 dig_ctrl_inst.latch_mem_inst.gclk\[9\] dig_ctrl_inst.latch_mem_inst.RAM\[9\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
X_1861_ VDPWR VGND VDPWR VGND _0523_ _0506_ _0278_ _0521_ _0463_ sky130_fd_sc_hd__o31ai_1
X_2413_ VGND VDPWR VDPWR VGND _1012_ dig_ctrl_inst.cpu_inst.port_o\[4\] net360 _0092_
+ sky130_fd_sc_hd__mux2_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[59\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[59\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[59\]._gclk sky130_fd_sc_hd__clkbuf_4
X_2344_ VGND VDPWR VDPWR VGND _0783_ net149 _0831_ _0983_ sky130_fd_sc_hd__o21ai_1
Xclkbuf_1_0__f_clk VGND VDPWR VDPWR VGND clknet_1_0__leaf_clk clknet_0_clk sky130_fd_sc_hd__clkbuf_16
X_1226_ VGND VDPWR VDPWR VGND net258 _1068_ _1035_ sky130_fd_sc_hd__nor2_1
X_2275_ VDPWR VGND VDPWR VGND dig_ctrl_inst.cpu_inst.data\[4\] _0916_ _0917_ _0813_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_59_150 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_5_Left_83 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2060_ VDPWR VGND VDPWR VGND net100 _0718_ dig_ctrl_inst.latch_mem_inst.RAM\[52\]\[7\]
+ net43 sky130_fd_sc_hd__and3_2
XFILLER_0_60_22 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
X_1913_ VDPWR VGND VDPWR VGND _0565_ _0278_ _0574_ _0556_ _0573_ sky130_fd_sc_hd__or4_1
X_1844_ VDPWR VGND VDPWR VGND _0500_ _0498_ _0506_ _0499_ _0505_ sky130_fd_sc_hd__or4_1
X_1775_ VGND VDPWR VDPWR VGND _0438_ net117 dig_ctrl_inst.latch_mem_inst.RAM\[49\]\[2\]
+ net138 net40 sky130_fd_sc_hd__and4_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[60\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND net178 dig_ctrl_inst.latch_mem_inst.gclk\[60\] dig_ctrl_inst.latch_mem_inst.RAM\[60\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
X_2258_ VDPWR VGND VDPWR VGND _0892_ _0901_ _0815_ _0893_ sky130_fd_sc_hd__and3_2
X_2327_ VGND VDPWR VDPWR VGND _0967_ _0953_ _0957_ _0819_ _0966_ sky130_fd_sc_hd__a211o_1
X_1209_ VDPWR VGND VDPWR VGND _1051_ dig_ctrl_inst.cpu_inst.rst_ni sky130_fd_sc_hd__inv_2
X_2189_ VGND VDPWR VDPWR VGND net149 _0798_ _0780_ _0834_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_153 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1560_ VDPWR VGND VDPWR VGND _0226_ dig_ctrl_inst.cpu_inst.regs\[1\]\[6\] _1035_
+ _1068_ dig_ctrl_inst.cpu_inst.regs\[2\]\[6\] _0225_ sky130_fd_sc_hd__a221o_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[30\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[30\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[30\]._gclk sky130_fd_sc_hd__clkbuf_4
X_1491_ VDPWR VGND VDPWR VGND _0178_ _0003_ net347 sky130_fd_sc_hd__xor2_1
X_2112_ VGND VDPWR VDPWR VGND _0762_ _0647_ dig_ctrl_inst.cpu_inst.data\[5\] _0040_
+ sky130_fd_sc_hd__mux2_1
X_2043_ VGND VDPWR VDPWR VGND _0699_ _0702_ _0701_ dig_ctrl_inst.latch_mem_inst.RAM\[27\]\[6\]
+ _0130_ _0700_ sky130_fd_sc_hd__a2111o_1
X_1827_ VGND VDPWR VDPWR VGND _0489_ net78 dig_ctrl_inst.latch_mem_inst.RAM\[30\]\[3\]
+ net115 net69 sky130_fd_sc_hd__and4_1
XFILLER_0_17_337 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_32_329 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
X_1758_ VGND VDPWR VDPWR VGND _0421_ net88 dig_ctrl_inst.latch_mem_inst.RAM\[41\]\[2\]
+ net116 net48 sky130_fd_sc_hd__and4_1
X_1689_ VDPWR VGND VDPWR VGND net113 _0353_ dig_ctrl_inst.latch_mem_inst.RAM\[18\]\[1\]
+ net62 sky130_fd_sc_hd__and3_2
XFILLER_0_20_80 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[53\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND net189 dig_ctrl_inst.latch_mem_inst.gclk\[53\] dig_ctrl_inst.latch_mem_inst.RAM\[53\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[42\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND net207 dig_ctrl_inst.latch_mem_inst.gclk\[42\] dig_ctrl_inst.latch_mem_inst.RAM\[42\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_35_145 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
Xdig_ctrl_inst.latch_mem_inst.gen_words\[31\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND net223 dig_ctrl_inst.latch_mem_inst.gclk\[31\] dig_ctrl_inst.latch_mem_inst.RAM\[31\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
X_1474_ VGND VDPWR VDPWR VGND net176 _0168_ _0166_ dig_ctrl_inst.cpu_inst.regs\[0\]\[6\]
+ _0167_ sky130_fd_sc_hd__o22a_2
Xfanout209 VGND VDPWR VDPWR VGND net210 net209 sky130_fd_sc_hd__clkbuf_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[20\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND net243 dig_ctrl_inst.latch_mem_inst.gclk\[20\] dig_ctrl_inst.latch_mem_inst.RAM\[20\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
X_1612_ VDPWR VGND VDPWR VGND _0274_ _0275_ _0273_ _0276_ _0277_ sky130_fd_sc_hd__or4_4
XFILLER_0_1_201 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2592_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.cpu_state\[2\] net156 _0106_
+ clknet_leaf_10_clk sky130_fd_sc_hd__dfrtp_1
X_1543_ VDPWR VGND VDPWR VGND _0211_ _1045_ _0197_ _0205_ _0023_ sky130_fd_sc_hd__a22oi_1
X_2026_ VDPWR VGND VDPWR VGND _0685_ _0140_ dig_ctrl_inst.latch_mem_inst.RAM\[30\]\[6\]
+ dig_ctrl_inst.latch_mem_inst.RAM\[37\]\[6\] _0132_ _0684_ sky130_fd_sc_hd__a221o_1
XFILLER_0_32_115 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[57\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND net181 dig_ctrl_inst.latch_mem_inst.gclk\[57\] dig_ctrl_inst.latch_mem_inst.RAM\[57\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[2\].gen_latches\[0\].p_latch VGND VDPWR VDPWR
+ VGND net240 dig_ctrl_inst.latch_mem_inst.gclk\[2\] dig_ctrl_inst.latch_mem_inst.RAM\[2\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[46\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND net198 dig_ctrl_inst.latch_mem_inst.gclk\[46\] dig_ctrl_inst.latch_mem_inst.RAM\[46\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
Xinput9 VGND VDPWR VDPWR VGND net9 ui_in[6] sky130_fd_sc_hd__clkbuf_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[35\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND net212 dig_ctrl_inst.latch_mem_inst.gclk\[35\] dig_ctrl_inst.latch_mem_inst.RAM\[35\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_36_35 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_39_270 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[24\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND net230 dig_ctrl_inst.latch_mem_inst.gclk\[24\] dig_ctrl_inst.latch_mem_inst.RAM\[24\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
X_2575_ VGND VDPWR VDPWR VGND net26 net173 _0089_ clknet_leaf_6_clk sky130_fd_sc_hd__dfrtp_1
X_1457_ VDPWR VGND VDPWR VGND net71 dig_ctrl_inst.latch_mem_inst.data_we\[60\] net142
+ net37 sky130_fd_sc_hd__and3_2
X_1526_ VGND VDPWR VDPWR VGND _0191_ net165 dig_ctrl_inst.cpu_inst.data\[0\] _0198_
+ sky130_fd_sc_hd__mux2_1
X_1388_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[23\] _0128_ net143
+ sky130_fd_sc_hd__and2_1
X_2009_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[48\]\[6\] _0151_ _0668_
+ dig_ctrl_inst.latch_mem_inst.RAM\[58\]\[6\] _0158_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_131 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[6\].gen_latches\[1\].p_latch VGND VDPWR VDPWR
+ VGND net233 dig_ctrl_inst.latch_mem_inst.gclk\[6\] dig_ctrl_inst.latch_mem_inst.RAM\[6\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[23\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[23\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[23\]._gclk sky130_fd_sc_hd__clkbuf_4
X_2360_ VGND VDPWR VDPWR VGND _0991_ _0995_ net323 _0056_ sky130_fd_sc_hd__mux2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[39\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND net207 dig_ctrl_inst.latch_mem_inst.gclk\[39\] dig_ctrl_inst.latch_mem_inst.RAM\[39\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
X_1311_ VDPWR VGND VDPWR VGND net159 _1153_ sky130_fd_sc_hd__inv_2
X_2291_ VDPWR VGND VDPWR VGND _0907_ _0234_ _0931_ _0932_ sky130_fd_sc_hd__a21o_1
X_1242_ VGND VDPWR VDPWR VGND _1084_ net262 dig_ctrl_inst.cpu_inst.regs\[2\]\[0\]
+ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_10_Right_10 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[28\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND net224 dig_ctrl_inst.latch_mem_inst.gclk\[28\] dig_ctrl_inst.latch_mem_inst.RAM\[28\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
XANTENNA_25 VGND VDPWR VDPWR VGND net80 sky130_fd_sc_hd__diode_2
XANTENNA_14 VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[52\] sky130_fd_sc_hd__diode_2
XFILLER_0_63_3 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[17\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND net242 dig_ctrl_inst.latch_mem_inst.gclk\[17\] dig_ctrl_inst.latch_mem_inst.RAM\[17\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
X_2558_ VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_data_o\[2\] net175 _0082_ clknet_leaf_9_clk
+ sky130_fd_sc_hd__dfrtp_1
X_2489_ VDPWR VGND VDPWR VGND dig_ctrl_inst.cpu_inst.port_o\[3\] clknet_leaf_6_clk
+ _0015_ sky130_fd_sc_hd__dfxtp_1
X_1509_ VGND VDPWR VDPWR VGND _0186_ _0189_ dig_ctrl_inst.cpu_inst.skip sky130_fd_sc_hd__nor2_2
XFILLER_0_65_313 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1860_ VGND VDPWR VDPWR VGND _0522_ _0506_ _0463_ _0278_ _0521_ sky130_fd_sc_hd__o31a_1
Xinput12 VGND VDPWR VDPWR VGND net12 uio_in[1] sky130_fd_sc_hd__clkbuf_1
X_1791_ VDPWR VGND VDPWR VGND net74 _0454_ dig_ctrl_inst.latch_mem_inst.RAM\[28\]\[2\]
+ net67 sky130_fd_sc_hd__and3_2
X_2412_ VGND VDPWR VDPWR VGND _1012_ dig_ctrl_inst.cpu_inst.port_o\[3\] net28 _0091_
+ sky130_fd_sc_hd__mux2_1
X_2343_ VDPWR VGND VDPWR VGND _0979_ _0982_ _0980_ _0981_ sky130_fd_sc_hd__or3_1
X_2274_ VGND VDPWR VDPWR VGND _0844_ _0235_ _0805_ _0916_ net163 sky130_fd_sc_hd__a2bb2o_1
X_1225_ VDPWR VGND VDPWR VGND _1062_ _1067_ _1064_ _1066_ sky130_fd_sc_hd__or3_1
XFILLER_0_59_162 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_17_clk VGND VDPWR VDPWR VGND clknet_leaf_17_clk clknet_1_0__leaf_clk
+ sky130_fd_sc_hd__clkbuf_8
X_1989_ VGND VDPWR VDPWR VGND _0270_ _0647_ net246 _0032_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_69 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_29_313 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_71_113 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[61\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND net223 dig_ctrl_inst.latch_mem_inst.gclk\[61\] dig_ctrl_inst.latch_mem_inst.RAM\[61\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
X_1843_ VDPWR VGND VDPWR VGND _0503_ _0501_ _0505_ _0502_ _0504_ sky130_fd_sc_hd__or4_1
X_1912_ VGND VDPWR VDPWR VGND _0571_ _0573_ _0572_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_6_clk VGND VDPWR VDPWR VGND clknet_leaf_6_clk clknet_1_1__leaf_clk sky130_fd_sc_hd__clkbuf_8
Xdig_ctrl_inst.latch_mem_inst.genblk1\[3\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[3\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[3\]._gclk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_12_268 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_1774_ VDPWR VGND VDPWR VGND net125 _0437_ dig_ctrl_inst.latch_mem_inst.RAM\[12\]\[2\]
+ net71 sky130_fd_sc_hd__and3_2
XFILLER_0_8_35 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1208_ VGND VDPWR VDPWR VGND net175 _1051_ net306 sky130_fd_sc_hd__nand2b_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[50\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND net242 dig_ctrl_inst.latch_mem_inst.gclk\[50\] dig_ctrl_inst.latch_mem_inst.RAM\[50\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_71_Left_149 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2257_ VGND VDPWR VDPWR VGND _0900_ _0894_ _0897_ _0764_ _0899_ sky130_fd_sc_hd__a211o_1
XFILLER_0_20_290 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2326_ VDPWR VGND VDPWR VGND _0966_ _1062_ _1057_ _0959_ _0965_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_47_165 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2188_ VGND VDPWR VDPWR VGND _0833_ _0832_ _1129_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_273 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_7_251 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_14_16 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.genblk1\[16\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[16\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[16\]._gclk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_39_57 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_1490_ VGND VDPWR VDPWR VGND _0179_ _0002_ _0178_ sky130_fd_sc_hd__nor2_1
Xhold1 VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.wdata\[4\] net283 sky130_fd_sc_hd__dlygate4sd3_1
X_2042_ VGND VDPWR VDPWR VGND _0701_ net79 dig_ctrl_inst.latch_mem_inst.RAM\[46\]\[6\]
+ net114 net55 sky130_fd_sc_hd__and4_1
X_2111_ VDPWR VGND VDPWR VGND _0576_ _0763_ _0039_ _0762_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_29_143 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_8_Right_8 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1826_ VGND VDPWR VDPWR VGND _0488_ net114 dig_ctrl_inst.latch_mem_inst.RAM\[14\]\[3\]
+ net127 net76 sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_39_Right_39 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1757_ VDPWR VGND VDPWR VGND _0414_ _0420_ _0415_ _0419_ sky130_fd_sc_hd__or3_1
X_1688_ VDPWR VGND VDPWR VGND net81 _0352_ dig_ctrl_inst.latch_mem_inst.RAM\[26\]\[1\]
+ net62 sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[54\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND net228 dig_ctrl_inst.latch_mem_inst.gclk\[54\] dig_ctrl_inst.latch_mem_inst.RAM\[54\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
X_2309_ VGND VDPWR VDPWR VGND _0949_ _0767_ _0948_ _0950_ _0768_ sky130_fd_sc_hd__a2bb2o_1
XPHY_EDGE_ROW_48_Right_48 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_43_190 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_57_Right_57 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_66_Right_66 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_25_37 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1611_ VGND VDPWR VDPWR VGND _1188_ _0276_ _1180_ net126 net97 _1190_ sky130_fd_sc_hd__a2111o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[31\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND net189 dig_ctrl_inst.latch_mem_inst.gclk\[31\] dig_ctrl_inst.latch_mem_inst.RAM\[31\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_75_Right_75 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2591_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.cpu_state\[1\] net156 _0105_
+ clknet_leaf_9_clk sky130_fd_sc_hd__dfrtp_4
X_1473_ VDPWR VGND VDPWR VGND net255 net251 _0167_ _1049_ sky130_fd_sc_hd__a21oi_1
X_1542_ VDPWR VGND VDPWR VGND _0186_ _0211_ _0209_ _0210_ sky130_fd_sc_hd__o21bai_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[20\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND net210 dig_ctrl_inst.latch_mem_inst.gclk\[20\] dig_ctrl_inst.latch_mem_inst.RAM\[20\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
X_2025_ VGND VDPWR VDPWR VGND _0684_ net120 dig_ctrl_inst.latch_mem_inst.RAM\[5\]\[6\]
+ net130 net101 sky130_fd_sc_hd__and4_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[58\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND net220 dig_ctrl_inst.latch_mem_inst.gclk\[58\] dig_ctrl_inst.latch_mem_inst.RAM\[58\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
X_1809_ VDPWR VGND VDPWR VGND net135 _0471_ dig_ctrl_inst.latch_mem_inst.RAM\[48\]\[3\]
+ net43 sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[47\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND net243 dig_ctrl_inst.latch_mem_inst.gclk\[47\] dig_ctrl_inst.latch_mem_inst.RAM\[47\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[2\].gen_latches\[4\].p_latch VGND VDPWR VDPWR
+ VGND net204 dig_ctrl_inst.latch_mem_inst.gclk\[2\] dig_ctrl_inst.latch_mem_inst.RAM\[2\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[35\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND net179 dig_ctrl_inst.latch_mem_inst.gclk\[35\] dig_ctrl_inst.latch_mem_inst.RAM\[35\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
X_2574_ VGND VDPWR VDPWR VGND net25 net173 _0088_ clknet_leaf_6_clk sky130_fd_sc_hd__dfrtp_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[14\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[14\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[14\]._gclk clknet_leaf_1_clk sky130_fd_sc_hd__dlclkp_1
XFILLER_0_6_338 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[24\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND net195 dig_ctrl_inst.latch_mem_inst.gclk\[24\] dig_ctrl_inst.latch_mem_inst.RAM\[24\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
X_1525_ VGND VDPWR VDPWR VGND _0197_ _0195_ _1075_ _0193_ _0196_ sky130_fd_sc_hd__and4_2
X_1387_ VGND VDPWR VDPWR VGND net107 net103 net68 _0128_ sky130_fd_sc_hd__and3_4
X_1456_ VDPWR VGND VDPWR VGND _0160_ net38 net71 sky130_fd_sc_hd__and2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[13\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND net213 dig_ctrl_inst.latch_mem_inst.gclk\[13\] dig_ctrl_inst.latch_mem_inst.RAM\[13\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
X_2008_ VDPWR VGND VDPWR VGND _0661_ _0667_ _0662_ _0666_ sky130_fd_sc_hd__or3_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[62\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[62\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[62\]._gclk sky130_fd_sc_hd__clkbuf_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[6\].gen_latches\[5\].p_latch VGND VDPWR VDPWR
+ VGND net201 dig_ctrl_inst.latch_mem_inst.gclk\[6\] dig_ctrl_inst.latch_mem_inst.RAM\[6\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_51_277 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1310_ VGND VDPWR VDPWR VGND _1061_ _1148_ _1149_ _1150_ _1151_ _1152_ sky130_fd_sc_hd__o41a_1
X_1241_ VDPWR VGND VDPWR VGND net258 _1083_ net262 dig_ctrl_inst.cpu_inst.regs\[3\]\[0\]
+ sky130_fd_sc_hd__and3_2
X_2290_ VGND VDPWR VDPWR VGND _0931_ _0930_ _0929_ sky130_fd_sc_hd__nand2_1
XANTENNA_15 VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_data_i\[2\] sky130_fd_sc_hd__diode_2
XANTENNA_26 VGND VDPWR VDPWR VGND net99 sky130_fd_sc_hd__diode_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[28\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND net190 dig_ctrl_inst.latch_mem_inst.gclk\[28\] dig_ctrl_inst.latch_mem_inst.RAM\[28\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
X_2557_ VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_data_o\[1\] net171 _0081_ clknet_leaf_5_clk
+ sky130_fd_sc_hd__dfrtp_1
X_1508_ VGND VDPWR VDPWR VGND _0188_ dig_ctrl_inst.cpu_inst.port_o\[7\] net324 _0011_
+ sky130_fd_sc_hd__mux2_1
X_2488_ VDPWR VGND VDPWR VGND dig_ctrl_inst.cpu_inst.port_o\[2\] clknet_leaf_6_clk
+ _0014_ sky130_fd_sc_hd__dfxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[17\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND net207 dig_ctrl_inst.latch_mem_inst.gclk\[17\] dig_ctrl_inst.latch_mem_inst.RAM\[17\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
X_1439_ VDPWR VGND VDPWR VGND net112 dig_ctrl_inst.latch_mem_inst.data_we\[50\] net143
+ net39 sky130_fd_sc_hd__and3_2
XFILLER_0_33_299 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_68_141 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xinput13 VGND VDPWR VDPWR VGND net13 uio_in[3] sky130_fd_sc_hd__clkbuf_1
X_1790_ VGND VDPWR VDPWR VGND _0453_ net79 dig_ctrl_inst.latch_mem_inst.RAM\[62\]\[2\]
+ net114 net45 sky130_fd_sc_hd__and4_1
X_2411_ VGND VDPWR VDPWR VGND _1012_ dig_ctrl_inst.cpu_inst.port_o\[2\] net27 _0090_
+ sky130_fd_sc_hd__mux2_1
X_1224_ VGND VDPWR VDPWR VGND _1066_ net258 net262 sky130_fd_sc_hd__nand2_1
X_2273_ VGND VDPWR VDPWR VGND _0914_ _0915_ _0913_ sky130_fd_sc_hd__nor2_1
X_2342_ VGND VDPWR VDPWR VGND _0975_ _0815_ _0764_ _0981_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_288 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1988_ VGND VDPWR VDPWR VGND _0648_ _0279_ _0578_ net33 sky130_fd_sc_hd__a21bo_1
X_2609_ VDPWR VGND VDPWR VGND uio_out[1] net273 sky130_fd_sc_hd__buf_2
XFILLER_0_65_100 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_0_119 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
Xfanout190 VGND VDPWR VDPWR VGND net191 net190 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_28_15 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_69 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1773_ VGND VDPWR VDPWR VGND _0433_ _0436_ _0435_ dig_ctrl_inst.latch_mem_inst.RAM\[33\]\[2\]
+ _0136_ _0434_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_44_339 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[61\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND net193 dig_ctrl_inst.latch_mem_inst.gclk\[61\] dig_ctrl_inst.latch_mem_inst.RAM\[61\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
X_1842_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[12\]\[3\] _0116_ _0504_
+ dig_ctrl_inst.latch_mem_inst.RAM\[27\]\[3\] _0130_ sky130_fd_sc_hd__a22o_1
X_1911_ VDPWR VGND VDPWR VGND _0568_ _0566_ _0572_ _0567_ _0570_ sky130_fd_sc_hd__or4_1
XFILLER_0_12_214 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_3 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_2187_ VGND VDPWR VDPWR VGND _0830_ _0832_ _0831_ _0776_ _0782_ sky130_fd_sc_hd__o22a_1
X_2256_ VDPWR VGND VDPWR VGND _0899_ _0844_ net158 net160 _0812_ _0898_ sky130_fd_sc_hd__a221o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[50\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND net205 dig_ctrl_inst.latch_mem_inst.gclk\[50\] dig_ctrl_inst.latch_mem_inst.RAM\[50\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
X_2325_ VDPWR VGND VDPWR VGND _0815_ _0964_ _0965_ _0959_ sky130_fd_sc_hd__a21oi_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[55\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[55\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[55\]._gclk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_53_169 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
Xdig_ctrl_inst.latch_mem_inst.genblk1\[19\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[19\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[19\]._gclk clknet_leaf_16_clk sky130_fd_sc_hd__dlclkp_1
Xhold2 VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.wdata\[6\] net284 sky130_fd_sc_hd__dlygate4sd3_1
X_2041_ VDPWR VGND VDPWR VGND net94 _0700_ dig_ctrl_inst.latch_mem_inst.RAM\[22\]\[6\]
+ net67 sky130_fd_sc_hd__and3_2
X_2110_ VGND VDPWR VDPWR VGND _0762_ _0763_ dig_ctrl_inst.cpu_inst.data\[4\] sky130_fd_sc_hd__nor2_1
XFILLER_0_44_114 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_17_306 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_1756_ VGND VDPWR VDPWR VGND _0416_ _0419_ _0418_ dig_ctrl_inst.latch_mem_inst.RAM\[27\]\[2\]
+ _0130_ _0417_ sky130_fd_sc_hd__a2111o_1
X_1825_ VGND VDPWR VDPWR VGND _0487_ net118 dig_ctrl_inst.latch_mem_inst.RAM\[49\]\[3\]
+ net138 net43 sky130_fd_sc_hd__and4_1
XFILLER_0_4_222 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_2308_ VDPWR VGND VDPWR VGND dig_ctrl_inst.spi_data_o\[5\] _0183_ _0949_ dig_ctrl_inst.synchronizer_port_i_inst\[5\].out
+ _0824_ sky130_fd_sc_hd__a22o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[54\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND net198 dig_ctrl_inst.latch_mem_inst.gclk\[54\] dig_ctrl_inst.latch_mem_inst.RAM\[54\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
X_1687_ VDPWR VGND VDPWR VGND net133 _0351_ dig_ctrl_inst.latch_mem_inst.RAM\[32\]\[1\]
+ net48 sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.genblk1\[21\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[21\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[21\]._gclk clknet_leaf_18_clk sky130_fd_sc_hd__dlclkp_1
X_2239_ VGND VDPWR VDPWR VGND _0772_ _0048_ _0876_ dig_ctrl_inst.cpu_inst.regs\[0\]\[2\]
+ _0882_ sky130_fd_sc_hd__o22a_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[43\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND net211 dig_ctrl_inst.latch_mem_inst.gclk\[43\] dig_ctrl_inst.latch_mem_inst.RAM\[43\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_35_169 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_8_3 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
Xdig_ctrl_inst.latch_mem_inst.gen_words\[32\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND net229 dig_ctrl_inst.latch_mem_inst.gclk\[32\] dig_ctrl_inst.latch_mem_inst.RAM\[32\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
X_2590_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.cpu_state\[0\] net153 _0104_
+ clknet_leaf_10_clk sky130_fd_sc_hd__dfrtp_4
X_1610_ VDPWR VGND VDPWR VGND _0117_ _0113_ _0275_ _0116_ _0118_ sky130_fd_sc_hd__or4_1
XFILLER_0_1_225 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1472_ VGND VDPWR VDPWR VGND net251 _0165_ net255 dig_ctrl_inst.cpu_inst.regs\[3\]\[6\]
+ _0166_ sky130_fd_sc_hd__a31o_1
XFILLER_0_1_247 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1541_ VGND VDPWR VDPWR VGND _0191_ net163 dig_ctrl_inst.cpu_inst.data\[3\] _0210_
+ sky130_fd_sc_hd__mux2_1
X_2024_ VGND VDPWR VDPWR VGND _0680_ _0683_ _0682_ dig_ctrl_inst.latch_mem_inst.RAM\[47\]\[6\]
+ _0149_ _0681_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_31_70 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_1808_ VGND VDPWR VDPWR VGND _0470_ net103 dig_ctrl_inst.latch_mem_inst.RAM\[21\]\[3\]
+ net117 net60 sky130_fd_sc_hd__and4_1
X_1739_ VDPWR VGND VDPWR VGND net97 _0402_ dig_ctrl_inst.latch_mem_inst.RAM\[52\]\[2\]
+ net41 sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[58\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND net187 dig_ctrl_inst.latch_mem_inst.gclk\[58\] dig_ctrl_inst.latch_mem_inst.RAM\[58\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[47\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND net209 dig_ctrl_inst.latch_mem_inst.gclk\[47\] dig_ctrl_inst.latch_mem_inst.RAM\[47\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[36\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND net226 dig_ctrl_inst.latch_mem_inst.gclk\[36\] dig_ctrl_inst.latch_mem_inst.RAM\[36\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[25\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND net236 dig_ctrl_inst.latch_mem_inst.gclk\[25\] dig_ctrl_inst.latch_mem_inst.RAM\[25\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_input_latches\[0\].n_latch VGND VDPWR VDPWR VGND
+ dig_ctrl_inst.data_out\[0\] clknet_leaf_9_clk dig_ctrl_inst.latch_mem_inst.wdata\[0\]
+ sky130_fd_sc_hd__dlxtn_1
XFILLER_0_54_220 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
X_1524_ VDPWR VGND VDPWR VGND _1036_ net245 _0196_ _1037_ sky130_fd_sc_hd__a21oi_1
X_2573_ VGND VDPWR VDPWR VGND dig_ctrl_inst.stb_d net175 dig_ctrl_inst.cpu_inst.stb_o
+ clknet_leaf_9_clk sky130_fd_sc_hd__dfrtp_1
X_1455_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[59\] _0159_ net147
+ sky130_fd_sc_hd__and2_1
X_1386_ VDPWR VGND VDPWR VGND net95 dig_ctrl_inst.latch_mem_inst.data_we\[22\] net145
+ net67 sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.genblk1\[48\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[48\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[48\]._gclk sky130_fd_sc_hd__clkbuf_4
X_2007_ VGND VDPWR VDPWR VGND _0663_ _0666_ _0665_ dig_ctrl_inst.latch_mem_inst.RAM\[9\]\[6\]
+ _1188_ _0664_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_45_220 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[13\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND net178 dig_ctrl_inst.latch_mem_inst.gclk\[13\] dig_ctrl_inst.latch_mem_inst.RAM\[13\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[7\].gen_latches\[0\].p_latch VGND VDPWR VDPWR
+ VGND net242 dig_ctrl_inst.latch_mem_inst.gclk\[7\] dig_ctrl_inst.latch_mem_inst.RAM\[7\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
X_1240_ VDPWR VGND VDPWR VGND _1037_ _1082_ _1036_ net245 sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[29\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND net230 dig_ctrl_inst.latch_mem_inst.gclk\[29\] dig_ctrl_inst.latch_mem_inst.RAM\[29\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
XANTENNA_16 VGND VDPWR VDPWR VGND net18 sky130_fd_sc_hd__diode_2
XANTENNA_27 VGND VDPWR VDPWR VGND net118 sky130_fd_sc_hd__diode_2
XFILLER_0_6_136 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2556_ VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_data_o\[0\] net171 _0080_ clknet_leaf_5_clk
+ sky130_fd_sc_hd__dfrtp_1
X_1507_ VGND VDPWR VDPWR VGND _0188_ dig_ctrl_inst.cpu_inst.port_o\[6\] net308 _0010_
+ sky130_fd_sc_hd__mux2_1
X_2487_ VDPWR VGND VDPWR VGND dig_ctrl_inst.cpu_inst.port_o\[1\] clknet_leaf_6_clk
+ _0013_ sky130_fd_sc_hd__dfxtp_1
X_1369_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[14\] _0118_ net145
+ sky130_fd_sc_hd__and2_1
X_1438_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[49\] _0152_ net148
+ sky130_fd_sc_hd__and2_1
Xinput14 VGND VDPWR VDPWR VGND net14 uio_in[4] sky130_fd_sc_hd__buf_1
X_2410_ VGND VDPWR VDPWR VGND _1012_ dig_ctrl_inst.cpu_inst.port_o\[1\] net26 _0089_
+ sky130_fd_sc_hd__mux2_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[3\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[3\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[3\]._gclk clknet_leaf_19_clk sky130_fd_sc_hd__dlclkp_1
X_2341_ VGND VDPWR VDPWR VGND _0980_ _0817_ _0976_ _0224_ _0978_ sky130_fd_sc_hd__a211o_1
X_2272_ VDPWR VGND VDPWR VGND _0914_ _0892_ net158 sky130_fd_sc_hd__and2_1
X_1223_ VGND VDPWR VDPWR VGND net176 _1065_ _1062_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_337 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.genblk1\[26\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[26\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[26\]._gclk clknet_leaf_19_clk sky130_fd_sc_hd__dlclkp_1
XFILLER_0_15_234 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_1987_ VDPWR VGND VDPWR VGND _0647_ _0279_ _0578_ net33 sky130_fd_sc_hd__a21boi_1
X_2608_ VDPWR VGND VDPWR VGND uio_out[0] net272 sky130_fd_sc_hd__buf_2
X_2539_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[2\]\[3\] net154 _0065_
+ clknet_leaf_12_clk sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_304 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xfanout180 VGND VDPWR VDPWR VGND net185 net180 sky130_fd_sc_hd__clkbuf_2
Xfanout191 VGND VDPWR VDPWR VGND net192 net191 sky130_fd_sc_hd__clkbuf_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[62\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND net228 dig_ctrl_inst.latch_mem_inst.gclk\[62\] dig_ctrl_inst.latch_mem_inst.RAM\[62\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
X_1910_ VDPWR VGND VDPWR VGND _0571_ _0143_ dig_ctrl_inst.latch_mem_inst.RAM\[13\]\[4\]
+ dig_ctrl_inst.latch_mem_inst.RAM\[40\]\[4\] _0117_ _0569_ sky130_fd_sc_hd__a221o_1
XFILLER_0_29_337 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1772_ VDPWR VGND VDPWR VGND net98 _0435_ dig_ctrl_inst.latch_mem_inst.RAM\[36\]\[2\]
+ net56 sky130_fd_sc_hd__and3_2
X_1841_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[3\]\[3\] _1180_ _0503_
+ dig_ctrl_inst.latch_mem_inst.RAM\[63\]\[3\] _0163_ sky130_fd_sc_hd__a22o_1
X_2324_ VDPWR VGND VDPWR VGND _0962_ _0960_ _0961_ _0964_ _0963_ sky130_fd_sc_hd__or4b_1
X_1206_ VDPWR VGND VDPWR VGND dig_ctrl_inst.port_ms_sync_i _1050_ sky130_fd_sc_hd__inv_2
X_2186_ VGND VDPWR VDPWR VGND _0831_ _0785_ net149 sky130_fd_sc_hd__nand2_1
X_2255_ VGND VDPWR VDPWR VGND _0806_ _0818_ _0898_ _1113_ _0241_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_34_81 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_9_Left_87 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xhold3 VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.wdata\[2\] net285 sky130_fd_sc_hd__dlygate4sd3_1
X_2040_ VDPWR VGND VDPWR VGND net86 _0699_ dig_ctrl_inst.latch_mem_inst.RAM\[56\]\[6\]
+ net45 sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[55\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND net236 dig_ctrl_inst.latch_mem_inst.gclk\[55\] dig_ctrl_inst.latch_mem_inst.RAM\[55\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
X_1824_ VDPWR VGND VDPWR VGND net98 _0486_ dig_ctrl_inst.latch_mem_inst.RAM\[36\]\[3\]
+ net56 sky130_fd_sc_hd__and3_2
X_1755_ VGND VDPWR VDPWR VGND _0418_ net76 dig_ctrl_inst.latch_mem_inst.RAM\[61\]\[2\]
+ net123 net43 sky130_fd_sc_hd__and4_1
X_1686_ VDPWR VGND VDPWR VGND _0348_ _0346_ _0350_ _0347_ _0349_ sky130_fd_sc_hd__or4_1
X_2307_ VGND VDPWR VDPWR VGND _0924_ _0948_ _1152_ sky130_fd_sc_hd__xnor2_1
X_2238_ VGND VDPWR VDPWR VGND _0882_ _0881_ _0880_ _0768_ _0771_ sky130_fd_sc_hd__a211o_1
X_2169_ VGND VDPWR VDPWR VGND _1076_ _0815_ _1060_ sky130_fd_sc_hd__nor2_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[43\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND net179 dig_ctrl_inst.latch_mem_inst.gclk\[43\] dig_ctrl_inst.latch_mem_inst.RAM\[43\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[32\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND net195 dig_ctrl_inst.latch_mem_inst.gclk\[32\] dig_ctrl_inst.latch_mem_inst.RAM\[32\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[21\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND net211 dig_ctrl_inst.latch_mem_inst.gclk\[21\] dig_ctrl_inst.latch_mem_inst.RAM\[21\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[12\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[12\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[12\]._gclk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_237 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
X_1540_ VDPWR VGND VDPWR VGND _0186_ _0209_ dig_ctrl_inst.cpu_inst.ip\[3\] _0204_
+ sky130_fd_sc_hd__and3_2
X_1471_ VGND VDPWR VDPWR VGND _0165_ net255 dig_ctrl_inst.cpu_inst.regs\[2\]\[6\]
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_66_68 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[59\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND net233 dig_ctrl_inst.latch_mem_inst.gclk\[59\] dig_ctrl_inst.latch_mem_inst.RAM\[59\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
X_2023_ VDPWR VGND VDPWR VGND net130 _0682_ dig_ctrl_inst.latch_mem_inst.RAM\[8\]\[6\]
+ net86 sky130_fd_sc_hd__and3_2
XPHY_EDGE_ROW_59_Left_137 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[10\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND net228 dig_ctrl_inst.latch_mem_inst.gclk\[10\] dig_ctrl_inst.latch_mem_inst.RAM\[10\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
X_1807_ VGND VDPWR VDPWR VGND _0469_ net88 dig_ctrl_inst.latch_mem_inst.RAM\[43\]\[3\]
+ net104 net50 sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_68_Left_146 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1669_ VGND VDPWR VDPWR VGND _0334_ net105 dig_ctrl_inst.latch_mem_inst.RAM\[15\]\[0\]
+ net132 net75 sky130_fd_sc_hd__and4_1
X_1738_ VDPWR VGND VDPWR VGND net133 _0401_ dig_ctrl_inst.latch_mem_inst.RAM\[32\]\[2\]
+ net52 sky130_fd_sc_hd__and3_2
XFILLER_0_0_281 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_181 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_77_Left_155 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[3\].gen_latches\[3\].p_latch VGND VDPWR VDPWR
+ VGND net212 dig_ctrl_inst.latch_mem_inst.gclk\[3\] dig_ctrl_inst.latch_mem_inst.RAM\[3\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[36\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND net190 dig_ctrl_inst.latch_mem_inst.gclk\[36\] dig_ctrl_inst.latch_mem_inst.RAM\[36\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[8\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[8\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[8\]._gclk clknet_leaf_0_clk sky130_fd_sc_hd__dlclkp_1
Xdig_ctrl_inst.latch_mem_inst.gen_input_latches\[4\].n_latch VDPWR VGND VDPWR VGND
+ dig_ctrl_inst.data_out\[4\] clknet_leaf_3_clk dig_ctrl_inst.latch_mem_inst.wdata\[4\]
+ sky130_fd_sc_hd__dlxtn_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[25\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND net203 dig_ctrl_inst.latch_mem_inst.gclk\[25\] dig_ctrl_inst.latch_mem_inst.RAM\[25\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_14_118 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2572_ VGND VDPWR VDPWR VGND dig_ctrl_inst.stb_dd net175 net304 clknet_leaf_9_clk
+ sky130_fd_sc_hd__dfrtp_1
X_1454_ VDPWR VGND VDPWR VGND net90 _0159_ net108 net46 sky130_fd_sc_hd__and3_2
X_1523_ VGND VDPWR VDPWR VGND _1072_ _0195_ _0194_ sky130_fd_sc_hd__or2_1
X_1385_ VDPWR VGND VDPWR VGND _0127_ net70 net93 sky130_fd_sc_hd__and2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[14\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND net219 dig_ctrl_inst.latch_mem_inst.gclk\[14\] dig_ctrl_inst.latch_mem_inst.RAM\[14\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
X_2006_ VDPWR VGND VDPWR VGND net84 _0665_ dig_ctrl_inst.latch_mem_inst.RAM\[24\]\[6\]
+ net60 sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.genblk1\[33\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[33\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[33\]._gclk clknet_leaf_4_clk sky130_fd_sc_hd__dlclkp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[7\].gen_latches\[4\].p_latch VGND VDPWR VDPWR
+ VGND net283 dig_ctrl_inst.latch_mem_inst.gclk\[7\] dig_ctrl_inst.latch_mem_inst.RAM\[7\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_36_221 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
Xdig_ctrl_inst.latch_mem_inst.gen_words\[29\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND net200 dig_ctrl_inst.latch_mem_inst.gclk\[29\] dig_ctrl_inst.latch_mem_inst.RAM\[29\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
XANTENNA_28 VGND VDPWR VDPWR VGND net227 sky130_fd_sc_hd__diode_2
XANTENNA_17 VGND VDPWR VDPWR VGND net103 sky130_fd_sc_hd__diode_2
XFILLER_0_27_221 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2555_ VDPWR VGND VDPWR VGND dig_ctrl_inst.spi_receiver_inst.stb_o clknet_leaf_5_clk
+ _0079_ sky130_fd_sc_hd__dfxtp_1
X_1506_ VGND VDPWR VDPWR VGND _0188_ dig_ctrl_inst.cpu_inst.port_o\[5\] net309 _0009_
+ sky130_fd_sc_hd__mux2_1
X_2486_ VDPWR VGND VDPWR VGND dig_ctrl_inst.cpu_inst.port_o\[0\] clknet_leaf_6_clk
+ _0012_ sky130_fd_sc_hd__dfxtp_1
X_1437_ VDPWR VGND VDPWR VGND net119 _0152_ net136 net43 sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[18\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND net213 dig_ctrl_inst.latch_mem_inst.gclk\[18\] dig_ctrl_inst.latch_mem_inst.RAM\[18\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
X_1299_ VDPWR VGND VDPWR VGND _1141_ _1139_ _1123_ _1107_ _1090_ _1052_ sky130_fd_sc_hd__o2111a_1
X_1368_ VDPWR VGND VDPWR VGND net115 _0118_ net130 net79 sky130_fd_sc_hd__and3_2
XFILLER_0_5_181 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_56_327 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_3_107 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2271_ VGND VDPWR VDPWR VGND _0892_ _0913_ net158 sky130_fd_sc_hd__nor2_1
X_2340_ VGND VDPWR VDPWR VGND _0805_ _0222_ _0977_ _0979_ sky130_fd_sc_hd__o21ai_1
X_1222_ VGND VDPWR VDPWR VGND net253 _1064_ net249 sky130_fd_sc_hd__or2_1
X_1986_ VGND VDPWR VDPWR VGND _0645_ _0641_ _0646_ _0631_ _0636_ sky130_fd_sc_hd__nor4_1
Xclkbuf_leaf_9_clk VGND VDPWR VDPWR VGND clknet_leaf_9_clk clknet_1_1__leaf_clk sky130_fd_sc_hd__clkbuf_8
X_2607_ VDPWR VGND VDPWR VGND uio_oe[7] net281 sky130_fd_sc_hd__buf_2
X_2469_ VGND VDPWR VDPWR VGND dig_ctrl_inst.synchronizer_port_i_inst\[3\].out net171
+ net298 clknet_leaf_5_clk sky130_fd_sc_hd__dfrtp_1
X_2538_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[2\]\[2\] net153 _0064_
+ clknet_leaf_12_clk sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_39 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xfanout170 VGND VDPWR VDPWR VGND net171 net170 sky130_fd_sc_hd__clkbuf_2
Xfanout192 VGND VDPWR VDPWR VGND net192 net193 sky130_fd_sc_hd__buf_1
Xfanout181 VGND VDPWR VDPWR VGND net184 net181 sky130_fd_sc_hd__clkbuf_2
X_1840_ VGND VDPWR VDPWR VGND _0464_ _0502_ _0476_ dig_ctrl_inst.latch_mem_inst.RAM\[32\]\[3\]
+ _0135_ _0472_ sky130_fd_sc_hd__a2111o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[62\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND net196 dig_ctrl_inst.latch_mem_inst.gclk\[62\] dig_ctrl_inst.latch_mem_inst.RAM\[62\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
X_1771_ VDPWR VGND VDPWR VGND net87 _0434_ dig_ctrl_inst.latch_mem_inst.RAM\[24\]\[2\]
+ net68 sky130_fd_sc_hd__and3_2
XPHY_EDGE_ROW_31_Left_109 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[51\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND net218 dig_ctrl_inst.latch_mem_inst.gclk\[51\] dig_ctrl_inst.latch_mem_inst.RAM\[51\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
X_2323_ VDPWR VGND VDPWR VGND _0221_ _0812_ _0963_ _0231_ _0817_ sky130_fd_sc_hd__a22o_1
X_2254_ VGND VDPWR VDPWR VGND _0897_ _0896_ _0895_ sky130_fd_sc_hd__nand2_1
X_1205_ VDPWR VGND VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[1\]\[6\] _1049_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_40_Left_118 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_47_113 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2185_ VGND VDPWR VDPWR VGND net150 _0783_ _0778_ _0830_ sky130_fd_sc_hd__mux2_1
X_1969_ VGND VDPWR VDPWR VGND _0579_ _0629_ _0592_ dig_ctrl_inst.latch_mem_inst.RAM\[14\]\[5\]
+ _0118_ _0590_ sky130_fd_sc_hd__a2111o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[40\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND net228 dig_ctrl_inst.latch_mem_inst.gclk\[40\] dig_ctrl_inst.latch_mem_inst.RAM\[40\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_35_308 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xhold4 VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.wdata\[0\] net286 sky130_fd_sc_hd__dlygate4sd3_1
X_1823_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[17\]\[3\] _0122_ _0485_
+ dig_ctrl_inst.latch_mem_inst.RAM\[59\]\[3\] _0159_ sky130_fd_sc_hd__a22o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[55\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND net207 dig_ctrl_inst.latch_mem_inst.gclk\[55\] dig_ctrl_inst.latch_mem_inst.RAM\[55\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
X_1754_ VDPWR VGND VDPWR VGND net132 _0417_ dig_ctrl_inst.latch_mem_inst.RAM\[6\]\[2\]
+ net96 sky130_fd_sc_hd__and3_2
Xmax_cap123 VGND VDPWR VDPWR VGND net123 _1174_ sky130_fd_sc_hd__buf_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[38\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[38\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[38\]._gclk clknet_leaf_19_clk sky130_fd_sc_hd__dlclkp_1
X_1685_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[39\]\[1\] _0142_ _0349_
+ dig_ctrl_inst.latch_mem_inst.RAM\[47\]\[1\] _0149_ sky130_fd_sc_hd__a22o_1
X_2237_ VDPWR VGND VDPWR VGND dig_ctrl_inst.spi_data_o\[2\] _0183_ _0881_ dig_ctrl_inst.synchronizer_port_i_inst\[2\].out
+ _0824_ sky130_fd_sc_hd__a22o_1
X_2306_ VDPWR VGND VDPWR VGND _0947_ _0924_ net159 sky130_fd_sc_hd__and2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[44\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND net224 dig_ctrl_inst.latch_mem_inst.gclk\[44\] dig_ctrl_inst.latch_mem_inst.RAM\[44\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_24_3 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_2099_ VGND VDPWR VDPWR VGND _0757_ net53 dig_ctrl_inst.latch_mem_inst.RAM\[53\]\[7\]
+ _0154_ dig_ctrl_inst.latch_mem_inst.RAM\[44\]\[7\] net72 sky130_fd_sc_hd__a32o_1
X_2168_ VDPWR VGND VDPWR VGND net164 _0812_ _0814_ dig_ctrl_inst.cpu_inst.data\[0\]
+ _0813_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_72 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_17_Right_17 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[33\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND net240 dig_ctrl_inst.latch_mem_inst.gclk\[33\] dig_ctrl_inst.latch_mem_inst.RAM\[33\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_26_Right_26 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.genblk1\[51\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[51\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[51\]._gclk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_25_29 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
Xdig_ctrl_inst.latch_mem_inst.genblk1\[40\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[40\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[40\]._gclk clknet_leaf_17_clk sky130_fd_sc_hd__dlclkp_1
XFILLER_0_41_39 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_26_149 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_35_Right_35 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1470_ VDPWR VGND VDPWR VGND net266 dig_ctrl_inst.spi_data_o\[5\] dig_ctrl_inst.data_out\[5\]
+ _0164_ _1147_ sky130_fd_sc_hd__a22o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[21\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND net181 dig_ctrl_inst.latch_mem_inst.gclk\[21\] dig_ctrl_inst.latch_mem_inst.RAM\[21\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_44_Right_44 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[59\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND net201 dig_ctrl_inst.latch_mem_inst.gclk\[59\] dig_ctrl_inst.latch_mem_inst.RAM\[59\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_53_Right_53 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2022_ VGND VDPWR VDPWR VGND _0681_ net90 dig_ctrl_inst.latch_mem_inst.RAM\[57\]\[6\]
+ net120 net47 sky130_fd_sc_hd__and4_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[10\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND net197 dig_ctrl_inst.latch_mem_inst.gclk\[10\] dig_ctrl_inst.latch_mem_inst.RAM\[10\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
X_1806_ VGND VDPWR VDPWR VGND _0468_ net80 dig_ctrl_inst.latch_mem_inst.RAM\[61\]\[3\]
+ net118 net43 sky130_fd_sc_hd__and4_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[48\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND net215 dig_ctrl_inst.latch_mem_inst.gclk\[48\] dig_ctrl_inst.latch_mem_inst.RAM\[48\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_62_Right_62 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_40_141 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1737_ VDPWR VGND VDPWR VGND net135 _0400_ dig_ctrl_inst.latch_mem_inst.RAM\[16\]\[2\]
+ net62 sky130_fd_sc_hd__and3_2
X_1599_ VGND VDPWR VDPWR VGND _0232_ _0257_ _0260_ _0264_ _0256_ _0265_ sky130_fd_sc_hd__o41a_1
XFILLER_0_0_293 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_1668_ VGND VDPWR VDPWR VGND _0330_ _0333_ _0332_ dig_ctrl_inst.latch_mem_inst.RAM\[1\]\[0\]
+ _1175_ _0331_ sky130_fd_sc_hd__a2111o_1
XPHY_EDGE_ROW_71_Right_71 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[3\].gen_latches\[7\].p_latch VGND VDPWR VDPWR
+ VGND net182 dig_ctrl_inst.latch_mem_inst.gclk\[3\] dig_ctrl_inst.latch_mem_inst.RAM\[3\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[37\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND net234 dig_ctrl_inst.latch_mem_inst.gclk\[37\] dig_ctrl_inst.latch_mem_inst.RAM\[37\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_12_Left_90 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2571_ VGND VDPWR VDPWR VGND dig_ctrl_inst.mode_d net171 net306 clknet_leaf_4_clk
+ sky130_fd_sc_hd__dfrtp_1
X_1522_ VGND VDPWR VDPWR VGND net167 dig_ctrl_inst.stb_dd dig_ctrl_inst.stb_d _0194_
+ sky130_fd_sc_hd__mux2_1
X_1453_ VDPWR VGND VDPWR VGND net83 dig_ctrl_inst.latch_mem_inst.data_we\[58\] net142
+ net37 sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[14\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND net193 dig_ctrl_inst.latch_mem_inst.gclk\[14\] dig_ctrl_inst.latch_mem_inst.RAM\[14\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
X_1384_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[21\] _0126_ net148
+ sky130_fd_sc_hd__and2_1
X_2005_ VGND VDPWR VDPWR VGND _0664_ net88 dig_ctrl_inst.latch_mem_inst.RAM\[25\]\[6\]
+ net117 net59 sky130_fd_sc_hd__and4_1
XANTENNA_29 VGND VDPWR VDPWR VGND net28 sky130_fd_sc_hd__diode_2
XANTENNA_18 VGND VDPWR VDPWR VGND net227 sky130_fd_sc_hd__diode_2
X_2554_ VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_miso_o net168 _0078_ clknet_leaf_4_clk
+ sky130_fd_sc_hd__dfrtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[18\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND net181 dig_ctrl_inst.latch_mem_inst.gclk\[18\] dig_ctrl_inst.latch_mem_inst.RAM\[18\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
X_2485_ VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_data_i\[7\] net172 _0011_ clknet_leaf_6_clk
+ sky130_fd_sc_hd__dfrtp_1
X_1505_ VGND VDPWR VDPWR VGND _0188_ dig_ctrl_inst.cpu_inst.port_o\[4\] net317 _0008_
+ sky130_fd_sc_hd__mux2_1
X_1436_ VDPWR VGND VDPWR VGND net143 dig_ctrl_inst.latch_mem_inst.data_we\[48\] net134
+ net39 sky130_fd_sc_hd__and3_2
X_1367_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[13\] _0117_ net141
+ sky130_fd_sc_hd__and2_1
X_1298_ VGND VDPWR VDPWR VGND _1138_ _1140_ _1122_ sky130_fd_sc_hd__nor2_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[44\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[44\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[44\]._gclk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_56_339 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2270_ VDPWR VGND VDPWR VGND _1129_ _0912_ _0796_ _0911_ _0909_ sky130_fd_sc_hd__o2bb2a_1
X_1221_ VGND VDPWR VDPWR VGND _1063_ net253 net249 sky130_fd_sc_hd__nor2_4
X_1985_ VDPWR VGND VDPWR VGND _0643_ _0627_ _0645_ _0642_ _0644_ sky130_fd_sc_hd__or4_1
X_2606_ VDPWR VGND VDPWR VGND uio_oe[6] net280 sky130_fd_sc_hd__buf_2
X_2537_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[2\]\[1\] net155 _0063_
+ clknet_leaf_12_clk sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_141 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2468_ VGND VDPWR VDPWR VGND dig_ctrl_inst.synchronizer_port_i_inst\[3\].pipe\[0\]
+ net169 net6 clknet_leaf_4_clk sky130_fd_sc_hd__dfrtp_1
X_2399_ VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_receiver_inst.spi_cnt\[2\] _1011_
+ net171 _0178_ _0079_ sky130_fd_sc_hd__a31o_1
X_1419_ VDPWR VGND VDPWR VGND net84 _0143_ net49 sky130_fd_sc_hd__and2_2
Xdig_ctrl_inst.latch_mem_inst.genblk1\[45\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[45\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[45\]._gclk clknet_leaf_0_clk sky130_fd_sc_hd__dlclkp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[63\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND net241 dig_ctrl_inst.latch_mem_inst.gclk\[63\] dig_ctrl_inst.latch_mem_inst.RAM\[63\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
Xfanout171 VDPWR VGND VDPWR VGND net171 dig_ctrl_inst.latch_mem_inst.rst_ni sky130_fd_sc_hd__buf_2
Xfanout193 VGND VDPWR VDPWR VGND net194 net193 sky130_fd_sc_hd__clkbuf_2
Xfanout182 VGND VDPWR VDPWR VGND net184 net182 sky130_fd_sc_hd__clkbuf_2
Xfanout160 VDPWR VGND VDPWR VGND net160 _1136_ sky130_fd_sc_hd__buf_2
X_1770_ VDPWR VGND VDPWR VGND net95 _0433_ dig_ctrl_inst.latch_mem_inst.RAM\[22\]\[2\]
+ net68 sky130_fd_sc_hd__and3_2
XFILLER_0_69_69 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1204_ VDPWR VGND VDPWR VGND dig_ctrl_inst.mode_d _1048_ sky130_fd_sc_hd__inv_2
X_2184_ VGND VDPWR VDPWR VGND _0771_ dig_ctrl_inst.cpu_inst.regs\[0\]\[0\] _0829_
+ _0046_ sky130_fd_sc_hd__mux2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[51\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND net182 dig_ctrl_inst.latch_mem_inst.gclk\[51\] dig_ctrl_inst.latch_mem_inst.RAM\[51\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_18_62 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2322_ VDPWR VGND VDPWR VGND dig_ctrl_inst.cpu_inst.data\[6\] _0813_ _0962_ net159
+ _0844_ sky130_fd_sc_hd__a22o_1
X_2253_ VDPWR VGND VDPWR VGND dig_ctrl_inst.cpu_inst.data\[3\] _0896_ _0813_ _0240_
+ _0805_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_62_128 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[40\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND net202 dig_ctrl_inst.latch_mem_inst.gclk\[40\] dig_ctrl_inst.latch_mem_inst.RAM\[40\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
X_1968_ VGND VDPWR VDPWR VGND _0593_ _0628_ _0599_ dig_ctrl_inst.latch_mem_inst.RAM\[53\]\[5\]
+ _0154_ _0595_ sky130_fd_sc_hd__a2111o_1
X_1899_ VDPWR VGND VDPWR VGND _0560_ _0156_ dig_ctrl_inst.latch_mem_inst.RAM\[34\]\[4\]
+ dig_ctrl_inst.latch_mem_inst.RAM\[56\]\[4\] _0137_ _0527_ sky130_fd_sc_hd__a221o_1
XFILLER_0_11_261 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xhold5 VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.wdata\[5\] net287 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_125 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_29_169 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1753_ VDPWR VGND VDPWR VGND net113 _0416_ dig_ctrl_inst.latch_mem_inst.RAM\[34\]\[2\]
+ net52 sky130_fd_sc_hd__and3_2
X_1822_ VDPWR VGND VDPWR VGND net72 _0484_ dig_ctrl_inst.latch_mem_inst.RAM\[44\]\[3\]
+ net52 sky130_fd_sc_hd__and3_2
X_1684_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[8\]\[1\] _1187_ _0348_
+ dig_ctrl_inst.latch_mem_inst.RAM\[42\]\[1\] _0145_ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_83 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_17_3 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2305_ VGND VDPWR VDPWR VGND _0932_ _0945_ _0819_ _0933_ _0946_ sky130_fd_sc_hd__a31o_1
X_2167_ VDPWR VGND VDPWR VGND net248 _1059_ _1058_ net246 _0813_ sky130_fd_sc_hd__o211a_2
X_2236_ VGND VDPWR VDPWR VGND _0879_ _0880_ _0767_ sky130_fd_sc_hd__nor2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[44\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND net189 dig_ctrl_inst.latch_mem_inst.gclk\[44\] dig_ctrl_inst.latch_mem_inst.RAM\[44\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
X_2098_ VDPWR VGND VDPWR VGND _0756_ _0157_ dig_ctrl_inst.latch_mem_inst.RAM\[38\]\[7\]
+ dig_ctrl_inst.latch_mem_inst.RAM\[57\]\[7\] _0141_ _0724_ sky130_fd_sc_hd__a221o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[0\].gen_latches\[1\].p_latch VGND VDPWR VDPWR
+ VGND net230 dig_ctrl_inst.latch_mem_inst.gclk\[0\] dig_ctrl_inst.latch_mem_inst.RAM\[0\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[37\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[37\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[37\]._gclk sky130_fd_sc_hd__clkbuf_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[33\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND net206 dig_ctrl_inst.latch_mem_inst.gclk\[33\] dig_ctrl_inst.latch_mem_inst.RAM\[33\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[22\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND net226 dig_ctrl_inst.latch_mem_inst.gclk\[22\] dig_ctrl_inst.latch_mem_inst.RAM\[22\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[11\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND net240 dig_ctrl_inst.latch_mem_inst.gclk\[11\] dig_ctrl_inst.latch_mem_inst.RAM\[11\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
X_2021_ VDPWR VGND VDPWR VGND net82 _0680_ dig_ctrl_inst.latch_mem_inst.RAM\[42\]\[6\]
+ net58 sky130_fd_sc_hd__and3_2
XFILLER_0_15_52 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1805_ VDPWR VGND VDPWR VGND net81 _0467_ dig_ctrl_inst.latch_mem_inst.RAM\[26\]\[3\]
+ net63 sky130_fd_sc_hd__and3_2
XFILLER_0_40_153 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_1736_ VGND VDPWR VDPWR VGND _0270_ _0399_ net257 _0028_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_175 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_1598_ VDPWR VGND VDPWR VGND net246 _0264_ _0236_ _0263_ _0251_ sky130_fd_sc_hd__or4bb_1
X_1667_ VGND VDPWR VDPWR VGND _0332_ net89 dig_ctrl_inst.latch_mem_inst.RAM\[43\]\[0\]
+ net105 net51 sky130_fd_sc_hd__and4_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[48\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND net178 dig_ctrl_inst.latch_mem_inst.gclk\[48\] dig_ctrl_inst.latch_mem_inst.RAM\[48\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
X_2219_ VGND VDPWR VDPWR VGND _1129_ _0808_ _0806_ _0863_ sky130_fd_sc_hd__mux2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[4\].gen_latches\[2\].p_latch VGND VDPWR VDPWR
+ VGND net219 dig_ctrl_inst.latch_mem_inst.gclk\[4\] dig_ctrl_inst.latch_mem_inst.RAM\[4\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_23_109 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[37\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND net198 dig_ctrl_inst.latch_mem_inst.gclk\[37\] dig_ctrl_inst.latch_mem_inst.RAM\[37\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_16_150 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_31_142 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_31_164 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_16_183 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_31_175 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_3 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
Xdig_ctrl_inst.latch_mem_inst.gen_words\[26\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND net215 dig_ctrl_inst.latch_mem_inst.gclk\[26\] dig_ctrl_inst.latch_mem_inst.RAM\[26\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
X_2570_ VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_receiver_inst.spi_sclk_sync net168
+ net297 clknet_leaf_4_clk sky130_fd_sc_hd__dfrtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[15\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND net234 dig_ctrl_inst.latch_mem_inst.gclk\[15\] dig_ctrl_inst.latch_mem_inst.RAM\[15\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
X_1383_ VDPWR VGND VDPWR VGND net102 _0126_ net119 net63 sky130_fd_sc_hd__and3_2
X_1521_ VGND VDPWR VDPWR VGND _0192_ dig_ctrl_inst.cpu_inst.skip _0185_ _0193_ sky130_fd_sc_hd__o21ai_1
X_1452_ VDPWR VGND VDPWR VGND _0158_ net39 net83 sky130_fd_sc_hd__and2_1
X_2004_ VGND VDPWR VDPWR VGND _0663_ net103 dig_ctrl_inst.latch_mem_inst.RAM\[21\]\[6\]
+ net117 net60 sky130_fd_sc_hd__and4_1
XFILLER_0_42_94 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_9_103 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
Xdig_ctrl_inst.latch_mem_inst.gen_words\[8\].gen_latches\[3\].p_latch VGND VDPWR VDPWR
+ VGND net215 dig_ctrl_inst.latch_mem_inst.gclk\[8\] dig_ctrl_inst.latch_mem_inst.RAM\[8\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
X_1719_ VDPWR VGND VDPWR VGND net98 _0383_ dig_ctrl_inst.latch_mem_inst.RAM\[52\]\[1\]
+ net46 sky130_fd_sc_hd__and3_2
XFILLER_0_36_278 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
Xdig_ctrl_inst.latch_mem_inst.genblk1\[52\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[52\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[52\]._gclk clknet_leaf_3_clk sky130_fd_sc_hd__dlclkp_1
XFILLER_0_59_337 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XANTENNA_19 VGND VDPWR VDPWR VGND net290 sky130_fd_sc_hd__diode_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[19\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND net223 dig_ctrl_inst.latch_mem_inst.gclk\[19\] dig_ctrl_inst.latch_mem_inst.RAM\[19\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
X_1504_ VGND VDPWR VDPWR VGND _0188_ dig_ctrl_inst.cpu_inst.port_o\[3\] dig_ctrl_inst.spi_data_i\[3\]
+ _0007_ sky130_fd_sc_hd__mux2_1
X_2553_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[3\]\[7\] net156 _0077_
+ clknet_leaf_8_clk sky130_fd_sc_hd__dfrtp_1
X_2484_ VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_data_i\[6\] net172 _0010_ clknet_leaf_5_clk
+ sky130_fd_sc_hd__dfrtp_1
X_1366_ VGND VDPWR VDPWR VGND net124 net116 net76 _0117_ sky130_fd_sc_hd__and3_4
X_1435_ VDPWR VGND VDPWR VGND _0151_ net39 net134 sky130_fd_sc_hd__and2_1
X_1297_ VGND VDPWR VDPWR VGND _1139_ _1137_ net264 _1043_ _1124_ _1131_ sky130_fd_sc_hd__a32o_1
X_2606__280 VGND VDPWR VDPWR VGND _2606__280/LO net280 sky130_fd_sc_hd__conb_1
X_1220_ VDPWR VGND VDPWR VGND net248 dig_ctrl_inst.cpu_inst.instr\[6\] net246 dig_ctrl_inst.cpu_inst.instr\[7\]
+ _1062_ sky130_fd_sc_hd__or4_4
XFILLER_0_23_52 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1984_ VGND VDPWR VDPWR VGND _0582_ _0644_ _0608_ dig_ctrl_inst.latch_mem_inst.RAM\[19\]\[5\]
+ _0124_ _0587_ sky130_fd_sc_hd__a2111o_1
X_2467_ VGND VDPWR VDPWR VGND dig_ctrl_inst.synchronizer_port_i_inst\[4\].out net169
+ net293 clknet_leaf_4_clk sky130_fd_sc_hd__dfrtp_1
X_2536_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[2\]\[0\] net156 _0062_
+ clknet_leaf_8_clk sky130_fd_sc_hd__dfrtp_1
X_2605_ VDPWR VGND VDPWR VGND uio_oe[5] net271 sky130_fd_sc_hd__buf_2
X_2398_ VGND VDPWR VDPWR VGND _1011_ net171 dig_ctrl_inst.spi_receiver_inst.stb_o
+ sky130_fd_sc_hd__and2b_1
X_1349_ VDPWR VGND VDPWR VGND net107 _1184_ net131 net103 sky130_fd_sc_hd__and3_2
X_1418_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[39\] _0142_ net145
+ sky130_fd_sc_hd__and2_1
XFILLER_0_3_51 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xfanout172 VGND VDPWR VDPWR VGND net172 net174 sky130_fd_sc_hd__clkbuf_4
Xfanout183 VGND VDPWR VDPWR VGND net183 net184 sky130_fd_sc_hd__buf_1
Xfanout150 VGND VDPWR VDPWR VGND net150 _1080_ sky130_fd_sc_hd__clkbuf_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[63\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND net206 dig_ctrl_inst.latch_mem_inst.gclk\[63\] dig_ctrl_inst.latch_mem_inst.RAM\[63\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
Xfanout194 VGND VDPWR VDPWR VGND net194 net284 sky130_fd_sc_hd__buf_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[52\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND net227 dig_ctrl_inst.latch_mem_inst.gclk\[52\] dig_ctrl_inst.latch_mem_inst.RAM\[52\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
X_2321_ VGND VDPWR VDPWR VGND _0805_ _0810_ _0961_ _0230_ _0229_ sky130_fd_sc_hd__o22ai_1
X_2183_ VGND VDPWR VDPWR VGND _0829_ _0828_ _0822_ sky130_fd_sc_hd__nand2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[41\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND net237 dig_ctrl_inst.latch_mem_inst.gclk\[41\] dig_ctrl_inst.latch_mem_inst.RAM\[41\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
X_2252_ VGND VDPWR VDPWR VGND _0808_ _0895_ _0810_ _1114_ _0239_ sky130_fd_sc_hd__o22a_1
X_1203_ VDPWR VGND VDPWR VGND dig_ctrl_inst.cpu_inst.ip\[5\] _1047_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_181 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_62_107 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1967_ VDPWR VGND VDPWR VGND _0620_ _0583_ _0627_ _0589_ _0625_ sky130_fd_sc_hd__or4_2
X_1898_ VGND VDPWR VDPWR VGND _0559_ _0133_ _0557_ dig_ctrl_inst.latch_mem_inst.RAM\[31\]\[4\]
+ _0558_ sky130_fd_sc_hd__a211o_1
X_2519_ VDPWR VGND VDPWR VGND dig_ctrl_inst.cpu_inst.prev_state\[2\] clknet_leaf_8_clk
+ _0045_ sky130_fd_sc_hd__dfxtp_1
Xhold6 VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.wdata\[7\] net288 sky130_fd_sc_hd__dlygate4sd3_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[56\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND net211 dig_ctrl_inst.latch_mem_inst.gclk\[56\] dig_ctrl_inst.latch_mem_inst.RAM\[56\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
X_1752_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[47\]\[2\] _0149_ _0415_
+ dig_ctrl_inst.latch_mem_inst.RAM\[53\]\[2\] _0154_ sky130_fd_sc_hd__a22o_1
X_1821_ VDPWR VGND VDPWR VGND net127 _0483_ dig_ctrl_inst.latch_mem_inst.RAM\[8\]\[3\]
+ net86 sky130_fd_sc_hd__and3_2
XFILLER_0_20_64 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_37_181 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_10_clk VGND VDPWR VDPWR VGND clknet_leaf_10_clk clknet_1_0__leaf_clk
+ sky130_fd_sc_hd__clkbuf_8
X_1683_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[13\]\[1\] _0117_ _0347_
+ dig_ctrl_inst.latch_mem_inst.RAM\[56\]\[1\] _0156_ sky130_fd_sc_hd__a22o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[45\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND net232 dig_ctrl_inst.latch_mem_inst.gclk\[45\] dig_ctrl_inst.latch_mem_inst.RAM\[45\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
X_2304_ VDPWR VGND VDPWR VGND _0940_ _0945_ _0941_ _0944_ sky130_fd_sc_hd__or3_1
X_2097_ VDPWR VGND VDPWR VGND _0753_ _0751_ _0755_ _0752_ _0754_ sky130_fd_sc_hd__or4_1
X_2166_ VGND VDPWR VDPWR VGND net249 net253 _1060_ _0812_ sky130_fd_sc_hd__nor3b_4
X_2235_ VGND VDPWR VDPWR VGND _0877_ _0879_ _0878_ sky130_fd_sc_hd__or2_1
XFILLER_0_16_321 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_3_Right_3 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[0\].gen_latches\[5\].p_latch VGND VDPWR VDPWR
+ VGND net198 dig_ctrl_inst.latch_mem_inst.gclk\[0\] dig_ctrl_inst.latch_mem_inst.RAM\[0\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_0_52 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_clk VGND VDPWR VDPWR VGND clknet_1_1__leaf_clk clknet_0_clk sky130_fd_sc_hd__clkbuf_16
Xdig_ctrl_inst.latch_mem_inst.genblk1\[57\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[57\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[57\]._gclk clknet_leaf_0_clk sky130_fd_sc_hd__dlclkp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[22\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND net191 dig_ctrl_inst.latch_mem_inst.gclk\[22\] dig_ctrl_inst.latch_mem_inst.RAM\[22\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
X_2020_ VGND VDPWR VDPWR VGND _0676_ _0679_ _0678_ dig_ctrl_inst.latch_mem_inst.RAM\[51\]\[6\]
+ _0153_ _0677_ sky130_fd_sc_hd__a2111o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[11\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND net207 dig_ctrl_inst.latch_mem_inst.gclk\[11\] dig_ctrl_inst.latch_mem_inst.RAM\[11\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_28_Left_106 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_40_187 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_40_165 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1804_ VDPWR VGND VDPWR VGND net84 _0466_ dig_ctrl_inst.latch_mem_inst.RAM\[56\]\[3\]
+ net38 sky130_fd_sc_hd__and3_2
X_1666_ VDPWR VGND VDPWR VGND net97 _0331_ dig_ctrl_inst.latch_mem_inst.RAM\[52\]\[0\]
+ net40 sky130_fd_sc_hd__and3_2
X_1735_ VDPWR VGND VDPWR VGND net34 _0399_ _0398_ _0279_ dig_ctrl_inst.latch_mem_inst.RAM\[0\]\[1\]
+ sky130_fd_sc_hd__o2bb2a_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[49\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND net219 dig_ctrl_inst.latch_mem_inst.gclk\[49\] dig_ctrl_inst.latch_mem_inst.RAM\[49\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_37_Left_115 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1597_ VGND VDPWR VDPWR VGND net164 _0263_ _1098_ sky130_fd_sc_hd__xnor2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[4\].gen_latches\[6\].p_latch VGND VDPWR VDPWR
+ VGND net193 dig_ctrl_inst.latch_mem_inst.gclk\[4\] dig_ctrl_inst.latch_mem_inst.RAM\[4\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[38\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND net237 dig_ctrl_inst.latch_mem_inst.gclk\[38\] dig_ctrl_inst.latch_mem_inst.RAM\[38\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
X_2149_ VDPWR VGND VDPWR VGND _0793_ _0795_ _1098_ sky130_fd_sc_hd__or2_2
X_2218_ VGND VDPWR VDPWR VGND _0786_ _0862_ _0776_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_46_Left_124 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_55_Left_133 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_31_187 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_64_Left_142 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[26\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND net182 dig_ctrl_inst.latch_mem_inst.gclk\[26\] dig_ctrl_inst.latch_mem_inst.RAM\[26\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_73_Left_151 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1520_ VDPWR VGND VDPWR VGND _1065_ _0191_ _0192_ _1068_ sky130_fd_sc_hd__a21oi_1
X_1382_ VDPWR VGND VDPWR VGND net98 dig_ctrl_inst.latch_mem_inst.data_we\[20\] net147
+ net68 sky130_fd_sc_hd__and3_2
X_1451_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[57\] _0157_ net145
+ sky130_fd_sc_hd__and2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[15\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND net196 dig_ctrl_inst.latch_mem_inst.gclk\[15\] dig_ctrl_inst.latch_mem_inst.RAM\[15\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_26_41 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2003_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[29\]\[6\] _0131_ _0662_
+ dig_ctrl_inst.latch_mem_inst.RAM\[60\]\[6\] _0160_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_268 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1718_ VDPWR VGND VDPWR VGND net129 _0382_ dig_ctrl_inst.latch_mem_inst.RAM\[6\]\[1\]
+ net94 sky130_fd_sc_hd__and3_2
X_1649_ VGND VDPWR VDPWR VGND _0311_ _0314_ _0313_ dig_ctrl_inst.latch_mem_inst.RAM\[17\]\[0\]
+ _0122_ _0312_ sky130_fd_sc_hd__a2111o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[8\].gen_latches\[7\].p_latch VGND VDPWR VDPWR
+ VGND net181 dig_ctrl_inst.latch_mem_inst.gclk\[8\] dig_ctrl_inst.latch_mem_inst.RAM\[8\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[19\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND net188 dig_ctrl_inst.latch_mem_inst.gclk\[19\] dig_ctrl_inst.latch_mem_inst.RAM\[19\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
X_2552_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[3\]\[6\] dig_ctrl_inst.cpu_inst.rst_ni
+ _0076_ clknet_leaf_5_clk sky130_fd_sc_hd__dfrtp_1
X_2483_ VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_data_i\[5\] net174 _0009_ clknet_leaf_5_clk
+ sky130_fd_sc_hd__dfrtp_1
X_1503_ VGND VDPWR VDPWR VGND _0188_ dig_ctrl_inst.cpu_inst.port_o\[2\] dig_ctrl_inst.spi_data_i\[2\]
+ _0006_ sky130_fd_sc_hd__mux2_1
X_1434_ VDPWR VGND VDPWR VGND _0150_ _1170_ _1156_ sky130_fd_sc_hd__and2_1
X_1296_ VGND VDPWR VDPWR VGND _1137_ _1131_ _1124_ _1043_ _1138_ net264 sky130_fd_sc_hd__a32oi_4
X_1365_ VDPWR VGND VDPWR VGND net148 dig_ctrl_inst.latch_mem_inst.data_we\[12\] net127
+ net73 sky130_fd_sc_hd__and3_2
XFILLER_0_5_151 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1207__1 VDPWR VGND VDPWR VGND clknet_leaf_5_clk net282 sky130_fd_sc_hd__inv_2
XFILLER_0_59_113 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2604_ VDPWR VGND VDPWR VGND uio_oe[4] net270 sky130_fd_sc_hd__buf_2
X_1983_ VGND VDPWR VDPWR VGND _0606_ _0643_ _0610_ dig_ctrl_inst.latch_mem_inst.RAM\[2\]\[5\]
+ _1178_ _0609_ sky130_fd_sc_hd__a2111o_1
X_2535_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[1\]\[7\] net156 _0061_
+ clknet_leaf_8_clk sky130_fd_sc_hd__dfrtp_1
X_2466_ VGND VDPWR VDPWR VGND dig_ctrl_inst.synchronizer_port_i_inst\[4\].pipe\[0\]
+ net170 net7 clknet_leaf_4_clk sky130_fd_sc_hd__dfrtp_1
X_1417_ VDPWR VGND VDPWR VGND net101 _0142_ net109 net58 sky130_fd_sc_hd__and3_2
X_2397_ VGND VDPWR VDPWR VGND _1004_ net330 _1010_ _0078_ sky130_fd_sc_hd__mux2_1
X_1279_ VGND VDPWR VDPWR VGND net264 _1120_ net167 _1121_ sky130_fd_sc_hd__a21oi_2
X_1348_ VDPWR VGND VDPWR VGND net143 dig_ctrl_inst.latch_mem_inst.data_we\[6\] net125
+ net93 sky130_fd_sc_hd__and3_2
Xfanout173 VGND VDPWR VDPWR VGND net173 net174 sky130_fd_sc_hd__clkbuf_4
Xfanout184 VDPWR VGND VDPWR VGND net184 net185 sky130_fd_sc_hd__buf_2
Xfanout195 VGND VDPWR VDPWR VGND net197 net195 sky130_fd_sc_hd__clkbuf_2
Xfanout151 VGND VDPWR VDPWR VGND net151 net152 sky130_fd_sc_hd__clkbuf_4
Xdig_ctrl_inst.latch_mem_inst.genblk1\[40\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[40\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[40\]._gclk sky130_fd_sc_hd__clkbuf_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[52\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND net192 dig_ctrl_inst.latch_mem_inst.gclk\[52\] dig_ctrl_inst.latch_mem_inst.RAM\[52\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
X_2251_ VGND VDPWR VDPWR VGND _0894_ _0893_ _0892_ sky130_fd_sc_hd__nand2_1
X_2320_ VGND VDPWR VDPWR VGND _0168_ _0808_ _0806_ _0960_ sky130_fd_sc_hd__mux2_1
X_2182_ VDPWR VGND VDPWR VGND _0768_ _0828_ _0827_ _0767_ net166 sky130_fd_sc_hd__o2bb2a_1
X_1202_ VDPWR VGND VDPWR VGND dig_ctrl_inst.cpu_inst.ip\[4\] _1046_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_97 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1966_ VDPWR VGND VDPWR VGND _0626_ _0153_ dig_ctrl_inst.latch_mem_inst.RAM\[17\]\[5\]
+ dig_ctrl_inst.latch_mem_inst.RAM\[51\]\[5\] _0122_ _0597_ sky130_fd_sc_hd__a221o_1
XFILLER_0_34_85 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
Xdig_ctrl_inst.latch_mem_inst.gen_words\[41\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND net204 dig_ctrl_inst.latch_mem_inst.gclk\[41\] dig_ctrl_inst.latch_mem_inst.RAM\[41\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[30\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND net224 dig_ctrl_inst.latch_mem_inst.gclk\[30\] dig_ctrl_inst.latch_mem_inst.RAM\[30\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
X_1897_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[2\]\[4\] _1178_ _0558_
+ dig_ctrl_inst.latch_mem_inst.RAM\[15\]\[4\] _0119_ sky130_fd_sc_hd__a22o_1
X_2449_ VGND VDPWR VDPWR VGND _1025_ _1030_ _1044_ _1027_ _0110_ sky130_fd_sc_hd__a31o_1
X_2518_ VDPWR VGND VDPWR VGND dig_ctrl_inst.cpu_inst.prev_state\[1\] clknet_leaf_9_clk
+ _0044_ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_296 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_6_290 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
Xhold7 VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.wdata\[3\] net289 sky130_fd_sc_hd__dlygate4sd3_1
X_1820_ VGND VDPWR VDPWR VGND _0482_ net76 dig_ctrl_inst.latch_mem_inst.RAM\[29\]\[3\]
+ net118 net62 sky130_fd_sc_hd__and4_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[56\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND net178 dig_ctrl_inst.latch_mem_inst.gclk\[56\] dig_ctrl_inst.latch_mem_inst.RAM\[56\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
X_1751_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[13\]\[2\] _0117_ _0414_
+ dig_ctrl_inst.latch_mem_inst.RAM\[21\]\[2\] _0126_ sky130_fd_sc_hd__a22o_1
X_1682_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[31\]\[1\] _0133_ _0346_
+ dig_ctrl_inst.latch_mem_inst.RAM\[38\]\[1\] _0141_ sky130_fd_sc_hd__a22o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[45\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND net199 dig_ctrl_inst.latch_mem_inst.gclk\[45\] dig_ctrl_inst.latch_mem_inst.RAM\[45\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_29_41 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_2303_ VGND VDPWR VDPWR VGND _0836_ _0944_ _0909_ _1114_ net162 _0943_ sky130_fd_sc_hd__o221a_1
X_2234_ VDPWR VGND VDPWR VGND net166 _1136_ _0878_ _1104_ sky130_fd_sc_hd__a21oi_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[1\].gen_latches\[0\].p_latch VGND VDPWR VDPWR
+ VGND net239 dig_ctrl_inst.latch_mem_inst.gclk\[1\] dig_ctrl_inst.latch_mem_inst.RAM\[1\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
X_2096_ VGND VDPWR VDPWR VGND _0754_ net41 dig_ctrl_inst.latch_mem_inst.RAM\[21\]\[7\]
+ _0126_ dig_ctrl_inst.latch_mem_inst.RAM\[54\]\[7\] net96 sky130_fd_sc_hd__a32o_1
X_2165_ VGND VDPWR VDPWR VGND _0805_ _0811_ _0810_ _0809_ _0258_ _0259_ sky130_fd_sc_hd__o221a_1
XFILLER_0_28_193 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[34\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND net214 dig_ctrl_inst.latch_mem_inst.gclk\[34\] dig_ctrl_inst.latch_mem_inst.RAM\[34\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
X_1949_ VDPWR VGND VDPWR VGND net85 _0609_ dig_ctrl_inst.latch_mem_inst.RAM\[24\]\[5\]
+ net59 sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[23\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND net234 dig_ctrl_inst.latch_mem_inst.gclk\[23\] dig_ctrl_inst.latch_mem_inst.RAM\[23\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_13_Right_13 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_25_152 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_1803_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[18\]\[3\] _0123_ _0465_
+ dig_ctrl_inst.latch_mem_inst.RAM\[40\]\[3\] _0143_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_308 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_22_Right_22 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1734_ VGND VDPWR VDPWR VGND _0397_ _0380_ _0277_ _0271_ _0398_ sky130_fd_sc_hd__o211a_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[5\].gen_latches\[1\].p_latch VGND VDPWR VDPWR
+ VGND net228 dig_ctrl_inst.latch_mem_inst.gclk\[5\] dig_ctrl_inst.latch_mem_inst.RAM\[5\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[49\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND net188 dig_ctrl_inst.latch_mem_inst.gclk\[49\] dig_ctrl_inst.latch_mem_inst.RAM\[49\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
X_1596_ VGND VDPWR VDPWR VGND _0262_ net164 _1098_ sky130_fd_sc_hd__nand2_1
X_1665_ VDPWR VGND VDPWR VGND net134 _0330_ dig_ctrl_inst.latch_mem_inst.RAM\[48\]\[0\]
+ net40 sky130_fd_sc_hd__and3_2
XFILLER_0_22_3 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2217_ VGND VDPWR VDPWR VGND _0797_ _0860_ _0861_ _0859_ sky130_fd_sc_hd__or3b_1
XPHY_EDGE_ROW_31_Right_31 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[38\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND net207 dig_ctrl_inst.latch_mem_inst.gclk\[38\] dig_ctrl_inst.latch_mem_inst.RAM\[38\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
X_2079_ VDPWR VGND VDPWR VGND _0735_ _0733_ _0737_ _0734_ _0736_ sky130_fd_sc_hd__or4_1
X_2148_ VGND VDPWR VDPWR VGND _0793_ _0794_ _1098_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_299 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_40_Right_40 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_31_133 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_16_141 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[27\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND net222 dig_ctrl_inst.latch_mem_inst.gclk\[27\] dig_ctrl_inst.latch_mem_inst.RAM\[27\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[33\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[33\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[33\]._gclk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_54_269 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
Xdig_ctrl_inst.latch_mem_inst.gen_words\[16\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND net237 dig_ctrl_inst.latch_mem_inst.gclk\[16\] dig_ctrl_inst.latch_mem_inst.RAM\[16\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
X_1450_ VDPWR VGND VDPWR VGND net90 _0157_ net120 net47 sky130_fd_sc_hd__and3_2
X_1381_ VDPWR VGND VDPWR VGND _0125_ net66 net99 sky130_fd_sc_hd__and2_1
X_2002_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[15\]\[6\] _0119_ _0661_
+ dig_ctrl_inst.latch_mem_inst.RAM\[23\]\[6\] _0128_ sky130_fd_sc_hd__a22o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[9\].gen_latches\[2\].p_latch VGND VDPWR VDPWR
+ VGND net221 dig_ctrl_inst.latch_mem_inst.gclk\[9\] dig_ctrl_inst.latch_mem_inst.RAM\[9\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
X_1648_ VDPWR VGND VDPWR VGND net128 _0313_ dig_ctrl_inst.latch_mem_inst.RAM\[2\]\[0\]
+ net113 sky130_fd_sc_hd__and3_2
X_1717_ VDPWR VGND VDPWR VGND net100 _0381_ dig_ctrl_inst.latch_mem_inst.RAM\[20\]\[1\]
+ net65 sky130_fd_sc_hd__and3_2
X_1579_ VGND VDPWR VDPWR VGND net160 _0245_ _1129_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_16_Left_94 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_12_11 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1502_ VGND VDPWR VDPWR VGND _0188_ dig_ctrl_inst.cpu_inst.port_o\[1\] net322 _0005_
+ sky130_fd_sc_hd__mux2_1
X_2482_ VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_data_i\[4\] net172 _0008_ clknet_leaf_5_clk
+ sky130_fd_sc_hd__dfrtp_1
X_2551_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[3\]\[5\] net157 _0075_
+ clknet_leaf_7_clk sky130_fd_sc_hd__dfrtp_1
X_1433_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[47\] _0149_ net145
+ sky130_fd_sc_hd__and2_1
X_1295_ VGND VDPWR VDPWR VGND net264 _1136_ net167 _1137_ sky130_fd_sc_hd__a21oi_2
X_1364_ VDPWR VGND VDPWR VGND _0116_ net72 net126 sky130_fd_sc_hd__and2_1
XFILLER_0_77_169 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_5_141 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[60\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND net224 dig_ctrl_inst.latch_mem_inst.gclk\[60\] dig_ctrl_inst.latch_mem_inst.RAM\[60\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_1_Left_79 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_59_169 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1982_ VGND VDPWR VDPWR VGND _0600_ _0642_ _0607_ dig_ctrl_inst.latch_mem_inst.RAM\[37\]\[5\]
+ _0140_ _0605_ sky130_fd_sc_hd__a2111o_1
X_2534_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[1\]\[6\] dig_ctrl_inst.cpu_inst.rst_ni
+ _0060_ clknet_leaf_5_clk sky130_fd_sc_hd__dfrtp_1
X_2603_ VDPWR VGND VDPWR VGND uio_oe[3] net269 sky130_fd_sc_hd__buf_2
X_2396_ VGND VDPWR VDPWR VGND _1005_ _1010_ _1007_ dig_ctrl_inst.spi_receiver_inst.spi_cnt\[2\]
+ _1009_ sky130_fd_sc_hd__o22a_1
X_2465_ VGND VDPWR VDPWR VGND dig_ctrl_inst.synchronizer_port_i_inst\[5\].out net169
+ net301 clknet_leaf_4_clk sky130_fd_sc_hd__dfrtp_1
X_1347_ VDPWR VGND VDPWR VGND _1183_ _1138_ _1123_ _1106_ _1090_ _1052_ sky130_fd_sc_hd__o2111a_1
X_1416_ VDPWR VGND VDPWR VGND net95 dig_ctrl_inst.latch_mem_inst.data_we\[38\] net146
+ net55 sky130_fd_sc_hd__and3_2
X_1278_ VGND VDPWR VDPWR VGND net177 _1116_ _1117_ _1118_ _1119_ _1120_ sky130_fd_sc_hd__o41a_2
Xfanout174 VGND VDPWR VDPWR VGND net174 dig_ctrl_inst.latch_mem_inst.rst_ni sky130_fd_sc_hd__clkbuf_4
Xfanout130 VDPWR VGND VDPWR VGND net130 net131 sky130_fd_sc_hd__buf_2
Xdig_ctrl_inst.latch_mem_inst.genblk1\[26\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[26\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[26\]._gclk sky130_fd_sc_hd__clkbuf_4
Xfanout185 VDPWR VGND VDPWR VGND net185 net288 sky130_fd_sc_hd__buf_2
Xfanout152 VGND VDPWR VDPWR VGND net152 net155 sky130_fd_sc_hd__clkbuf_4
Xfanout163 VDPWR VGND VDPWR VGND net163 _1120_ sky130_fd_sc_hd__buf_2
Xfanout196 VGND VDPWR VDPWR VGND net197 net196 sky130_fd_sc_hd__clkbuf_2
Xfanout141 VGND VDPWR VDPWR VGND net142 net141 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_69_Right_69 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[53\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND net231 dig_ctrl_inst.latch_mem_inst.gclk\[53\] dig_ctrl_inst.latch_mem_inst.RAM\[53\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
X_2250_ VGND VDPWR VDPWR VGND _0893_ _0868_ net163 sky130_fd_sc_hd__nand2_1
X_1201_ VDPWR VGND VDPWR VGND dig_ctrl_inst.cpu_inst.ip\[3\] _1045_ sky130_fd_sc_hd__inv_2
X_2181_ VDPWR VGND VDPWR VGND _0827_ _0824_ dig_ctrl_inst.spi_data_o\[0\] dig_ctrl_inst.synchronizer_port_i_inst\[0\].out
+ _0183_ _0826_ sky130_fd_sc_hd__a221o_1
X_1965_ VDPWR VGND VDPWR VGND net74 _0625_ dig_ctrl_inst.latch_mem_inst.RAM\[28\]\[5\]
+ net66 sky130_fd_sc_hd__and3_2
XFILLER_0_34_97 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2517_ VDPWR VGND VDPWR VGND dig_ctrl_inst.cpu_inst.prev_state\[0\] clknet_leaf_8_clk
+ _0043_ sky130_fd_sc_hd__dfxtp_1
X_1896_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[12\]\[4\] _0116_ _0557_
+ dig_ctrl_inst.latch_mem_inst.RAM\[25\]\[4\] _0129_ sky130_fd_sc_hd__a22o_1
X_2379_ VGND VDPWR VDPWR VGND _1002_ _0999_ net338 _0068_ sky130_fd_sc_hd__mux2_1
X_2448_ VDPWR VGND VDPWR VGND _1030_ _1028_ dig_ctrl_inst.spi_addr\[3\] sky130_fd_sc_hd__and2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[30\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND net190 dig_ctrl_inst.latch_mem_inst.gclk\[30\] dig_ctrl_inst.latch_mem_inst.RAM\[30\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
Xhold8 VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.wdata\[1\] net290 sky130_fd_sc_hd__dlygate4sd3_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[57\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND net219 dig_ctrl_inst.latch_mem_inst.gclk\[57\] dig_ctrl_inst.latch_mem_inst.RAM\[57\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[46\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND net242 dig_ctrl_inst.latch_mem_inst.gclk\[46\] dig_ctrl_inst.latch_mem_inst.RAM\[46\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_37_150 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1750_ VDPWR VGND VDPWR VGND _0410_ _0413_ _0411_ _0412_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_4_Left_82 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1681_ VDPWR VGND VDPWR VGND _0343_ _0341_ _0345_ _0342_ _0344_ sky130_fd_sc_hd__or4_1
X_2233_ VDPWR VGND VDPWR VGND _1104_ _0877_ net166 _1136_ sky130_fd_sc_hd__and3_2
XFILLER_0_29_53 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.genblk1\[10\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[10\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[10\]._gclk clknet_leaf_17_clk sky130_fd_sc_hd__dlclkp_1
X_2164_ VGND VDPWR VDPWR VGND net246 net247 _0804_ _0810_ sky130_fd_sc_hd__or3b_4
X_2302_ VGND VDPWR VDPWR VGND _0883_ _0943_ _0942_ _0832_ _0857_ _0795_ sky130_fd_sc_hd__o221ai_1
X_2095_ VGND VDPWR VDPWR VGND _0753_ net63 dig_ctrl_inst.latch_mem_inst.RAM\[20\]\[7\]
+ _0125_ dig_ctrl_inst.latch_mem_inst.RAM\[26\]\[7\] net81 sky130_fd_sc_hd__a32o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[1\].gen_latches\[4\].p_latch VGND VDPWR VDPWR
+ VGND net208 dig_ctrl_inst.latch_mem_inst.gclk\[1\] dig_ctrl_inst.latch_mem_inst.RAM\[1\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_9_63 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
X_1879_ VDPWR VGND VDPWR VGND net85 _0540_ dig_ctrl_inst.latch_mem_inst.RAM\[24\]\[4\]
+ net59 sky130_fd_sc_hd__and3_2
XFILLER_0_31_315 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1948_ VGND VDPWR VDPWR VGND _0608_ net89 dig_ctrl_inst.latch_mem_inst.RAM\[25\]\[5\]
+ net117 net59 sky130_fd_sc_hd__and4_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[34\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND net178 dig_ctrl_inst.latch_mem_inst.gclk\[34\] dig_ctrl_inst.latch_mem_inst.RAM\[34\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_31_337 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[23\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND net201 dig_ctrl_inst.latch_mem_inst.gclk\[23\] dig_ctrl_inst.latch_mem_inst.RAM\[23\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[12\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND net212 dig_ctrl_inst.latch_mem_inst.gclk\[12\] dig_ctrl_inst.latch_mem_inst.RAM\[12\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_22_337 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_66_18 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1802_ VDPWR VGND VDPWR VGND net112 _0464_ dig_ctrl_inst.latch_mem_inst.RAM\[34\]\[3\]
+ net51 sky130_fd_sc_hd__and3_2
X_1733_ VGND VDPWR VDPWR VGND _0396_ _0392_ _0397_ _0384_ _0388_ sky130_fd_sc_hd__nor4_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[6\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[6\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[6\]._gclk sky130_fd_sc_hd__clkbuf_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[5\].gen_latches\[5\].p_latch VGND VDPWR VDPWR
+ VGND net202 dig_ctrl_inst.latch_mem_inst.gclk\[5\] dig_ctrl_inst.latch_mem_inst.RAM\[5\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
X_1595_ VGND VDPWR VDPWR VGND _1098_ _0261_ net164 sky130_fd_sc_hd__or2_1
XFILLER_0_13_337 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1664_ VGND VDPWR VDPWR VGND _0326_ _0329_ _0328_ dig_ctrl_inst.latch_mem_inst.RAM\[33\]\[0\]
+ _0136_ _0327_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_0_253 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_2216_ VGND VDPWR VDPWR VGND _0782_ _0860_ _0800_ _0781_ _0776_ sky130_fd_sc_hd__o22a_1
X_2147_ VDPWR VGND VDPWR VGND _1039_ _0793_ net247 _0774_ sky130_fd_sc_hd__or3_1
X_2078_ VGND VDPWR VDPWR VGND _0725_ _0736_ _0727_ dig_ctrl_inst.latch_mem_inst.RAM\[14\]\[7\]
+ _0118_ _0726_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_8_320 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_16_197 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.genblk1\[19\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[19\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[19\]._gclk sky130_fd_sc_hd__clkbuf_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[27\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND net191 dig_ctrl_inst.latch_mem_inst.gclk\[27\] dig_ctrl_inst.latch_mem_inst.RAM\[27\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[16\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND net208 dig_ctrl_inst.latch_mem_inst.gclk\[16\] dig_ctrl_inst.latch_mem_inst.RAM\[16\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_22_167 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1380_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[19\] _0124_ net141
+ sky130_fd_sc_hd__and2_1
X_2001_ VDPWR VGND VDPWR VGND _0658_ _0656_ _0660_ _0657_ _0659_ sky130_fd_sc_hd__or4_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[9\].gen_latches\[6\].p_latch VGND VDPWR VDPWR
+ VGND net186 dig_ctrl_inst.latch_mem_inst.gclk\[9\] dig_ctrl_inst.latch_mem_inst.RAM\[9\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
X_1716_ VGND VDPWR VDPWR VGND _0379_ _0375_ _0380_ _0369_ _0373_ sky130_fd_sc_hd__nor4_1
X_1647_ VDPWR VGND VDPWR VGND net94 _0312_ dig_ctrl_inst.latch_mem_inst.RAM\[22\]\[0\]
+ net65 sky130_fd_sc_hd__and3_2
X_1578_ VGND VDPWR VDPWR VGND _0244_ net160 _1129_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_3 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_59_318 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2550_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[3\]\[4\] net157 _0074_
+ clknet_leaf_7_clk sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_281 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
X_2481_ VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_data_i\[3\] net174 _0007_ clknet_leaf_5_clk
+ sky130_fd_sc_hd__dfrtp_1
X_1501_ VGND VDPWR VDPWR VGND _0188_ dig_ctrl_inst.cpu_inst.port_o\[0\] net337 _0004_
+ sky130_fd_sc_hd__mux2_1
X_1363_ VGND VDPWR VDPWR VGND _1138_ _1122_ _1090_ _1052_ _1107_ _0115_ sky130_fd_sc_hd__o2111a_2
XFILLER_0_50_262 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_1432_ VDPWR VGND VDPWR VGND net79 _0149_ net109 net58 sky130_fd_sc_hd__and3_2
XFILLER_0_37_97 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
X_1294_ VGND VDPWR VDPWR VGND net177 _1133_ _1134_ _1135_ _1132_ _1136_ sky130_fd_sc_hd__o41a_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[60\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND net188 dig_ctrl_inst.latch_mem_inst.gclk\[60\] dig_ctrl_inst.latch_mem_inst.RAM\[60\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_68_137 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.genblk1\[15\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[15\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[15\]._gclk clknet_leaf_15_clk sky130_fd_sc_hd__dlclkp_1
X_2613__276 VGND VDPWR VDPWR VGND net276 _2613__276/HI sky130_fd_sc_hd__conb_1
XFILLER_0_23_11 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1981_ VDPWR VGND VDPWR VGND _0639_ _0637_ _0641_ _0638_ _0640_ sky130_fd_sc_hd__or4_1
X_2533_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[1\]\[5\] net157 _0059_
+ clknet_leaf_7_clk sky130_fd_sc_hd__dfrtp_1
X_2602_ VDPWR VGND VDPWR VGND uio_oe[2] net279 sky130_fd_sc_hd__buf_2
XFILLER_0_2_178 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2395_ VGND VDPWR VDPWR VGND _1009_ dig_ctrl_inst.spi_receiver_inst.spi_cnt\[1\]
+ dig_ctrl_inst.spi_receiver_inst.spi_cnt\[2\] _1008_ sky130_fd_sc_hd__a21bo_1
X_2464_ VGND VDPWR VDPWR VGND dig_ctrl_inst.synchronizer_port_i_inst\[5\].pipe\[0\]
+ net170 net8 clknet_leaf_4_clk sky130_fd_sc_hd__dfrtp_1
X_1346_ VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[5\] net120 net130
+ net145 net101 sky130_fd_sc_hd__and4_1
X_1415_ VDPWR VGND VDPWR VGND _0141_ net53 net94 sky130_fd_sc_hd__and2_1
Xwire33 VGND VDPWR VDPWR VGND net33 _0646_ sky130_fd_sc_hd__clkbuf_1
X_1277_ VDPWR VGND VDPWR VGND net261 _1119_ net257 dig_ctrl_inst.cpu_inst.regs\[0\]\[3\]
+ sky130_fd_sc_hd__or3_1
XFILLER_0_14_240 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xfanout131 VGND VDPWR VDPWR VGND net132 net131 sky130_fd_sc_hd__clkbuf_2
Xfanout120 VGND VDPWR VDPWR VGND net122 net120 sky130_fd_sc_hd__clkbuf_2
Xfanout175 VGND VDPWR VDPWR VGND net175 dig_ctrl_inst.latch_mem_inst.rst_ni sky130_fd_sc_hd__clkbuf_4
Xfanout153 VGND VDPWR VDPWR VGND net153 net155 sky130_fd_sc_hd__clkbuf_4
Xfanout164 VGND VDPWR VDPWR VGND net164 _1104_ sky130_fd_sc_hd__clkbuf_4
Xfanout197 VGND VDPWR VDPWR VGND net198 net197 sky130_fd_sc_hd__clkbuf_2
Xfanout186 VGND VDPWR VDPWR VGND net187 net186 sky130_fd_sc_hd__clkbuf_2
Xfanout142 VDPWR VGND VDPWR VGND net144 net142 sky130_fd_sc_hd__dlymetal6s2s_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[53\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND net202 dig_ctrl_inst.latch_mem_inst.gclk\[53\] dig_ctrl_inst.latch_mem_inst.RAM\[53\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_37_310 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_69_29 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1200_ VDPWR VGND VDPWR VGND dig_ctrl_inst.spi_addr\[3\] _1044_ sky130_fd_sc_hd__inv_2
X_2180_ VGND VDPWR VDPWR VGND _0825_ _0826_ _1050_ sky130_fd_sc_hd__nor2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[42\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND net216 dig_ctrl_inst.latch_mem_inst.gclk\[42\] dig_ctrl_inst.latch_mem_inst.RAM\[42\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_47_129 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_1895_ VDPWR VGND VDPWR VGND _0550_ _0543_ _0556_ _0548_ _0555_ sky130_fd_sc_hd__or4_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[31\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND net231 dig_ctrl_inst.latch_mem_inst.gclk\[31\] dig_ctrl_inst.latch_mem_inst.RAM\[31\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
X_1964_ VDPWR VGND VDPWR VGND net124 _0624_ dig_ctrl_inst.latch_mem_inst.RAM\[12\]\[5\]
+ net71 sky130_fd_sc_hd__and3_2
Xclkbuf_leaf_13_clk VGND VDPWR VDPWR VGND clknet_leaf_13_clk clknet_1_0__leaf_clk
+ sky130_fd_sc_hd__clkbuf_8
X_2447_ VDPWR VGND VDPWR VGND _0109_ _1029_ _1028_ sky130_fd_sc_hd__and2_1
XFILLER_0_59_95 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2516_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.data\[7\] net151 _0042_ clknet_leaf_14_clk
+ sky130_fd_sc_hd__dfrtp_1
X_1329_ VGND VDPWR VDPWR VGND _1170_ _1171_ _1156_ sky130_fd_sc_hd__nor2_1
X_2378_ VGND VDPWR VDPWR VGND _1002_ _0998_ net321 _0067_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_107 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_46_173 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
Xhold9 VGND VDPWR VDPWR VGND dig_ctrl_inst.synchronizer_port_i_inst\[6\].pipe\[0\]
+ net291 sky130_fd_sc_hd__dlygate4sd3_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[57\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND net191 dig_ctrl_inst.latch_mem_inst.gclk\[57\] dig_ctrl_inst.latch_mem_inst.RAM\[57\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_29_107 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xmax_cap139 VDPWR VGND VDPWR VGND net139 _1013_ sky130_fd_sc_hd__buf_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[46\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND net208 dig_ctrl_inst.latch_mem_inst.gclk\[46\] dig_ctrl_inst.latch_mem_inst.RAM\[46\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
X_1680_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[40\]\[1\] _0143_ _0344_
+ dig_ctrl_inst.latch_mem_inst.RAM\[5\]\[1\] _0272_ sky130_fd_sc_hd__a22o_1
X_2301_ VGND VDPWR VDPWR VGND _1080_ _0780_ _0778_ _0942_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_2_clk VGND VDPWR VDPWR VGND clknet_leaf_2_clk clknet_1_1__leaf_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_29_65 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2163_ VGND VDPWR VDPWR VGND net150 _0808_ _0806_ _0809_ sky130_fd_sc_hd__mux2_1
X_2232_ VDPWR VGND VDPWR VGND _0871_ _0867_ _0876_ _0875_ _0874_ sky130_fd_sc_hd__or4b_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[35\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND net225 dig_ctrl_inst.latch_mem_inst.gclk\[35\] dig_ctrl_inst.latch_mem_inst.RAM\[35\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
X_2094_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[31\]\[7\] _0133_ _0752_
+ dig_ctrl_inst.latch_mem_inst.RAM\[55\]\[7\] _0155_ sky130_fd_sc_hd__a22o_1
X_1878_ VDPWR VGND VDPWR VGND net133 _0539_ dig_ctrl_inst.latch_mem_inst.RAM\[48\]\[4\]
+ net41 sky130_fd_sc_hd__and3_2
X_1947_ VGND VDPWR VDPWR VGND _0607_ net118 dig_ctrl_inst.latch_mem_inst.RAM\[49\]\[5\]
+ net138 net41 sky130_fd_sc_hd__and4_1
XFILLER_0_28_162 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[24\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND net243 dig_ctrl_inst.latch_mem_inst.gclk\[24\] dig_ctrl_inst.latch_mem_inst.RAM\[24\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[12\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND net182 dig_ctrl_inst.latch_mem_inst.gclk\[12\] dig_ctrl_inst.latch_mem_inst.RAM\[12\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
X_1732_ VGND VDPWR VDPWR VGND _0393_ _0396_ _0395_ dig_ctrl_inst.latch_mem_inst.RAM\[1\]\[1\]
+ _1175_ _0394_ sky130_fd_sc_hd__a2111o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[6\].gen_latches\[0\].p_latch VGND VDPWR VDPWR
+ VGND net240 dig_ctrl_inst.latch_mem_inst.gclk\[6\] dig_ctrl_inst.latch_mem_inst.RAM\[6\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_40_135 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_13_327 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_1801_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[0\]\[3\] _0463_ _0271_
+ _0277_ sky130_fd_sc_hd__or3_1
X_1663_ VGND VDPWR VDPWR VGND _0328_ net118 dig_ctrl_inst.latch_mem_inst.RAM\[13\]\[0\]
+ net126 net75 sky130_fd_sc_hd__and4_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[39\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND net218 dig_ctrl_inst.latch_mem_inst.gclk\[39\] dig_ctrl_inst.latch_mem_inst.RAM\[39\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
X_1594_ VGND VDPWR VDPWR VGND _0260_ _0258_ _0259_ sky130_fd_sc_hd__and2b_1
XFILLER_0_0_265 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Right_7 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2215_ VGND VDPWR VDPWR VGND net150 _0858_ _0788_ _0857_ _0859_ _0795_ sky130_fd_sc_hd__o32ai_2
X_2146_ VGND VDPWR VDPWR VGND _0791_ _0792_ _0789_ sky130_fd_sc_hd__nor2_1
X_2077_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[15\]\[7\] _0119_ _0735_
+ dig_ctrl_inst.latch_mem_inst.RAM\[23\]\[7\] _0128_ sky130_fd_sc_hd__a22o_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[58\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[58\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[58\]._gclk sky130_fd_sc_hd__clkbuf_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[28\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND net232 dig_ctrl_inst.latch_mem_inst.gclk\[28\] dig_ctrl_inst.latch_mem_inst.RAM\[28\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_31_113 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_2600__267 VGND VDPWR VDPWR VGND net267 _2600__267/HI sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_24_Left_102 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_33_Left_111 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_42_Left_120 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2000_ VGND VDPWR VDPWR VGND _0659_ net54 dig_ctrl_inst.latch_mem_inst.RAM\[16\]\[6\]
+ _0121_ dig_ctrl_inst.latch_mem_inst.RAM\[44\]\[6\] net72 sky130_fd_sc_hd__a32o_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[22\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[22\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[22\]._gclk clknet_leaf_0_clk sky130_fd_sc_hd__dlclkp_1
X_1646_ VGND VDPWR VDPWR VGND _0311_ net77 dig_ctrl_inst.latch_mem_inst.RAM\[45\]\[0\]
+ net122 net54 sky130_fd_sc_hd__and4_1
X_1715_ VGND VDPWR VDPWR VGND _0376_ _0379_ _0378_ dig_ctrl_inst.latch_mem_inst.RAM\[34\]\[1\]
+ _0137_ _0377_ sky130_fd_sc_hd__a2111o_1
X_1577_ VGND VDPWR VDPWR VGND _1099_ _0243_ net164 sky130_fd_sc_hd__or2_1
X_2129_ VGND VDPWR VDPWR VGND _0773_ _0775_ _0774_ sky130_fd_sc_hd__or2_1
X_2480_ VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_data_i\[2\] net174 _0006_ clknet_leaf_5_clk
+ sky130_fd_sc_hd__dfrtp_1
X_1500_ VGND VDPWR VDPWR VGND _0188_ _0184_ _0187_ sky130_fd_sc_hd__nor2_4
X_1362_ VGND VDPWR VDPWR VGND _1139_ _0114_ _1123_ sky130_fd_sc_hd__nor2_1
X_1431_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[46\] _0148_ net148
+ sky130_fd_sc_hd__and2_1
X_1293_ VGND VDPWR VDPWR VGND _1135_ net260 dig_ctrl_inst.cpu_inst.regs\[1\]\[2\]
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_53_53 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_33_219 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[61\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND net233 dig_ctrl_inst.latch_mem_inst.gclk\[61\] dig_ctrl_inst.latch_mem_inst.RAM\[61\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
X_1629_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[25\]\[0\] _0129_ _0294_
+ dig_ctrl_inst.latch_mem_inst.RAM\[62\]\[0\] _0162_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_165 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_23_78 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_1980_ VGND VDPWR VDPWR VGND _0585_ _0640_ _0598_ dig_ctrl_inst.latch_mem_inst.RAM\[13\]\[5\]
+ _0117_ _0586_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_23_23 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_2532_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[1\]\[4\] net157 _0058_
+ clknet_leaf_6_clk sky130_fd_sc_hd__dfrtp_1
X_2463_ VGND VDPWR VDPWR VGND dig_ctrl_inst.synchronizer_port_i_inst\[6\].out net169
+ net291 clknet_leaf_5_clk sky130_fd_sc_hd__dfrtp_1
X_2601_ VDPWR VGND VDPWR VGND uio_oe[1] net268 sky130_fd_sc_hd__buf_2
XFILLER_0_2_135 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2394_ VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_receiver_inst.spi_cnt\[0\] dig_ctrl_inst.spi_data_i\[0\]
+ dig_ctrl_inst.spi_data_i\[1\] _1008_ sky130_fd_sc_hd__mux2_1
X_1414_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[37\] _0140_ net145
+ sky130_fd_sc_hd__and2_1
X_1345_ VDPWR VGND VDPWR VGND net147 dig_ctrl_inst.latch_mem_inst.data_we\[4\] net129
+ net98 sky130_fd_sc_hd__and3_2
XFILLER_0_48_97 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1276_ VGND VDPWR VDPWR VGND _1118_ net257 dig_ctrl_inst.cpu_inst.regs\[1\]\[3\]
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_3_33 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_3_11 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_58_193 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xwire34 VGND VDPWR VDPWR VGND net34 _0365_ sky130_fd_sc_hd__clkbuf_1
Xfanout110 VGND VDPWR VDPWR VGND _1179_ net110 sky130_fd_sc_hd__clkbuf_2
Xfanout132 VGND VDPWR VDPWR VGND _1171_ net132 sky130_fd_sc_hd__clkbuf_2
Xfanout121 VGND VDPWR VDPWR VGND net122 net121 sky130_fd_sc_hd__clkbuf_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[54\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND net238 dig_ctrl_inst.latch_mem_inst.gclk\[54\] dig_ctrl_inst.latch_mem_inst.RAM\[54\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
Xfanout143 VGND VDPWR VDPWR VGND net144 net143 sky130_fd_sc_hd__clkbuf_2
Xfanout165 VGND VDPWR VDPWR VGND net165 _1087_ sky130_fd_sc_hd__clkbuf_4
Xfanout154 VGND VDPWR VDPWR VGND net155 net154 sky130_fd_sc_hd__clkbuf_2
Xfanout187 VGND VDPWR VDPWR VGND net187 net188 sky130_fd_sc_hd__buf_1
Xfanout198 VGND VDPWR VDPWR VGND net287 net198 sky130_fd_sc_hd__clkbuf_2
Xfanout176 VDPWR VGND VDPWR VGND net176 _1064_ sky130_fd_sc_hd__buf_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[42\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND net181 dig_ctrl_inst.latch_mem_inst.gclk\[42\] dig_ctrl_inst.latch_mem_inst.RAM\[42\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[31\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND net202 dig_ctrl_inst.latch_mem_inst.gclk\[31\] dig_ctrl_inst.latch_mem_inst.RAM\[31\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
X_1894_ VDPWR VGND VDPWR VGND _0553_ _0551_ _0555_ _0552_ _0554_ sky130_fd_sc_hd__or4_1
X_1963_ VDPWR VGND VDPWR VGND net133 _0623_ dig_ctrl_inst.latch_mem_inst.RAM\[16\]\[5\]
+ net61 sky130_fd_sc_hd__and3_2
X_2446_ VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_addr\[1\] dig_ctrl_inst.spi_addr\[2\]
+ dig_ctrl_inst.spi_addr\[0\] _1023_ _1029_ sky130_fd_sc_hd__a31o_1
X_2515_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.data\[6\] net151 _0041_ clknet_leaf_13_clk
+ sky130_fd_sc_hd__dfrtp_1
X_2377_ VGND VDPWR VDPWR VGND _1002_ _0997_ net331 _0066_ sky130_fd_sc_hd__mux2_1
X_1328_ VDPWR VGND VDPWR VGND _1170_ _1169_ _1157_ _1163_ dig_ctrl_inst.spi_addr\[4\]
+ _1041_ sky130_fd_sc_hd__o32a_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[20\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND net217 dig_ctrl_inst.latch_mem_inst.gclk\[20\] dig_ctrl_inst.latch_mem_inst.RAM\[20\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
X_1259_ VGND VDPWR VDPWR VGND _1101_ net257 dig_ctrl_inst.cpu_inst.regs\[1\]\[1\]
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_19_322 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[58\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND net230 dig_ctrl_inst.latch_mem_inst.gclk\[58\] dig_ctrl_inst.latch_mem_inst.RAM\[58\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[4\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[4\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[4\]._gclk clknet_leaf_4_clk sky130_fd_sc_hd__dlclkp_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[27\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[27\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[27\]._gclk clknet_leaf_1_clk sky130_fd_sc_hd__dlclkp_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[22\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[22\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[22\]._gclk sky130_fd_sc_hd__clkbuf_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[2\].gen_latches\[3\].p_latch VGND VDPWR VDPWR
+ VGND net212 dig_ctrl_inst.latch_mem_inst.gclk\[2\] dig_ctrl_inst.latch_mem_inst.RAM\[2\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
X_2231_ VGND VDPWR VDPWR VGND _1114_ _0861_ _0862_ net161 _0875_ sky130_fd_sc_hd__o211a_1
X_2300_ VGND VDPWR VDPWR VGND _0935_ _0815_ _0764_ _0941_ sky130_fd_sc_hd__mux2_1
X_2093_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[29\]\[7\] _0131_ _0751_
+ dig_ctrl_inst.latch_mem_inst.RAM\[62\]\[7\] _0162_ sky130_fd_sc_hd__a22o_1
X_2162_ VGND VDPWR VDPWR VGND net246 net247 _0808_ _0774_ sky130_fd_sc_hd__or3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[35\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND net189 dig_ctrl_inst.latch_mem_inst.gclk\[35\] dig_ctrl_inst.latch_mem_inst.RAM\[35\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_28_141 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1877_ VDPWR VGND VDPWR VGND net111 _0538_ dig_ctrl_inst.latch_mem_inst.RAM\[50\]\[4\]
+ net39 sky130_fd_sc_hd__and3_2
X_1946_ VDPWR VGND VDPWR VGND net125 _0606_ dig_ctrl_inst.latch_mem_inst.RAM\[4\]\[5\]
+ net97 sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[24\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND net205 dig_ctrl_inst.latch_mem_inst.gclk\[24\] dig_ctrl_inst.latch_mem_inst.RAM\[24\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
X_2429_ VGND VDPWR VDPWR VGND _0709_ _1017_ _1054_ _0462_ _0648_ _0761_ sky130_fd_sc_hd__a2111o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[13\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND net222 dig_ctrl_inst.latch_mem_inst.gclk\[13\] dig_ctrl_inst.latch_mem_inst.RAM\[13\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_57_225 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_15_57 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1800_ VGND VDPWR VDPWR VGND _0270_ _0462_ net253 _0029_ sky130_fd_sc_hd__mux2_1
X_1662_ VGND VDPWR VDPWR VGND _0327_ net105 dig_ctrl_inst.latch_mem_inst.RAM\[11\]\[0\]
+ net126 net92 sky130_fd_sc_hd__and4_1
X_1731_ VGND VDPWR VDPWR VGND _0395_ net90 dig_ctrl_inst.latch_mem_inst.RAM\[43\]\[1\]
+ net110 net54 sky130_fd_sc_hd__and4_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[6\].gen_latches\[4\].p_latch VGND VDPWR VDPWR
+ VGND net205 dig_ctrl_inst.latch_mem_inst.gclk\[6\] dig_ctrl_inst.latch_mem_inst.RAM\[6\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_0_277 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1593_ VGND VDPWR VDPWR VGND _0259_ net165 net150 sky130_fd_sc_hd__nand2_1
X_2214_ VGND VDPWR VDPWR VGND _0791_ net150 _0858_ _0799_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_48_203 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[39\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND net183 dig_ctrl_inst.latch_mem_inst.gclk\[39\] dig_ctrl_inst.latch_mem_inst.RAM\[39\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_72_63 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2076_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[9\]\[7\] _1188_ _0734_
+ dig_ctrl_inst.latch_mem_inst.RAM\[60\]\[7\] _0160_ sky130_fd_sc_hd__a22o_1
X_2145_ VGND VDPWR VDPWR VGND _0790_ _0791_ net149 sky130_fd_sc_hd__nor2_1
X_1929_ VDPWR VGND VDPWR VGND net95 _0589_ dig_ctrl_inst.latch_mem_inst.RAM\[22\]\[5\]
+ net67 sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[28\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND net199 dig_ctrl_inst.latch_mem_inst.gclk\[28\] dig_ctrl_inst.latch_mem_inst.RAM\[28\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_31_125 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
Xdig_ctrl_inst.latch_mem_inst.gen_words\[17\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND net217 dig_ctrl_inst.latch_mem_inst.gclk\[17\] dig_ctrl_inst.latch_mem_inst.RAM\[17\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_10_309 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_26_23 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_42_22 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
X_1645_ VGND VDPWR VDPWR VGND _0307_ _0310_ _0309_ dig_ctrl_inst.latch_mem_inst.RAM\[51\]\[0\]
+ _0153_ _0308_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_53_261 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_1576_ VGND VDPWR VDPWR VGND _0242_ net164 net149 _1099_ net165 sky130_fd_sc_hd__a211o_1
X_1714_ VDPWR VGND VDPWR VGND net97 _0378_ dig_ctrl_inst.latch_mem_inst.RAM\[36\]\[1\]
+ net50 sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.genblk1\[2\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[2\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[2\]._gclk sky130_fd_sc_hd__clkbuf_4
X_2059_ VDPWR VGND VDPWR VGND net127 _0717_ dig_ctrl_inst.latch_mem_inst.RAM\[12\]\[7\]
+ net73 sky130_fd_sc_hd__and3_2
X_2128_ VGND VDPWR VDPWR VGND _0774_ dig_ctrl_inst.cpu_inst.instr\[6\] dig_ctrl_inst.cpu_inst.instr\[7\]
+ sky130_fd_sc_hd__nand2b_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[15\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[15\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[15\]._gclk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_50_242 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_1430_ VDPWR VGND VDPWR VGND net75 _0148_ net114 net52 sky130_fd_sc_hd__and3_2
XFILLER_0_2_328 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_1361_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[11\] _0113_ net148
+ sky130_fd_sc_hd__and2_1
XFILLER_0_37_77 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1292_ VGND VDPWR VDPWR VGND net263 net260 _1134_ dig_ctrl_inst.cpu_inst.regs\[2\]\[2\]
+ sky130_fd_sc_hd__and3b_1
X_1559_ VDPWR VGND VDPWR VGND net258 _0225_ net262 dig_ctrl_inst.cpu_inst.regs\[3\]\[6\]
+ sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[61\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND net201 dig_ctrl_inst.latch_mem_inst.gclk\[61\] dig_ctrl_inst.latch_mem_inst.RAM\[61\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_68_3 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1628_ VDPWR VGND VDPWR VGND _0290_ _0293_ _0291_ _0292_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_61_Left_139 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.genblk1\[9\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[9\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[9\]._gclk clknet_leaf_16_clk sky130_fd_sc_hd__dlclkp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[50\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND net211 dig_ctrl_inst.latch_mem_inst.gclk\[50\] dig_ctrl_inst.latch_mem_inst.RAM\[50\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_70_Left_148 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_17_294 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_35 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2600_ VDPWR VGND VDPWR VGND uio_oe[0] net267 sky130_fd_sc_hd__buf_2
XFILLER_0_23_57 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_23_68 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2393_ VGND VDPWR VDPWR VGND _1007_ dig_ctrl_inst.spi_receiver_inst.spi_cnt\[1\]
+ _1006_ sky130_fd_sc_hd__and2b_1
X_2462_ VGND VDPWR VDPWR VGND dig_ctrl_inst.synchronizer_port_i_inst\[6\].pipe\[0\]
+ net168 net9 clknet_leaf_4_clk sky130_fd_sc_hd__dfrtp_1
X_1413_ VDPWR VGND VDPWR VGND net101 _0140_ net121 net56 sky130_fd_sc_hd__and3_2
X_2531_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[1\]\[3\] net154 _0057_
+ clknet_leaf_12_clk sky130_fd_sc_hd__dfrtp_1
X_1344_ VDPWR VGND VDPWR VGND _1182_ _1138_ _1123_ _1107_ _1090_ _1052_ sky130_fd_sc_hd__o2111a_1
Xwire35 VGND VDPWR VDPWR VGND net35 _0707_ sky130_fd_sc_hd__clkbuf_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[34\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[34\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[34\]._gclk clknet_leaf_16_clk sky130_fd_sc_hd__dlclkp_1
X_1275_ VGND VDPWR VDPWR VGND _1117_ net261 dig_ctrl_inst.cpu_inst.regs\[2\]\[3\]
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_61_337 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xfanout144 VGND VDPWR VDPWR VGND _1173_ net144 sky130_fd_sc_hd__clkbuf_2
Xfanout122 VGND VDPWR VDPWR VGND _1174_ net122 sky130_fd_sc_hd__clkbuf_2
Xfanout100 VGND VDPWR VDPWR VGND _1182_ net100 sky130_fd_sc_hd__clkbuf_2
Xfanout166 VDPWR VGND VDPWR VGND _1087_ net166 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout199 VGND VDPWR VDPWR VGND net200 net199 sky130_fd_sc_hd__clkbuf_2
Xfanout188 VDPWR VGND VDPWR VGND net188 net189 sky130_fd_sc_hd__buf_2
Xfanout111 VDPWR VGND VDPWR VGND net111 net113 sky130_fd_sc_hd__buf_2
Xfanout133 VDPWR VGND VDPWR VGND net133 net135 sky130_fd_sc_hd__buf_2
Xfanout155 VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.rst_ni net155 sky130_fd_sc_hd__clkbuf_2
Xfanout177 VDPWR VGND VDPWR VGND net177 _1061_ sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_29_Right_29 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[54\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND net205 dig_ctrl_inst.latch_mem_inst.gclk\[54\] dig_ctrl_inst.latch_mem_inst.RAM\[54\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_38_Right_38 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[43\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND net219 dig_ctrl_inst.latch_mem_inst.gclk\[43\] dig_ctrl_inst.latch_mem_inst.RAM\[43\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_47_Right_47 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[32\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND net238 dig_ctrl_inst.latch_mem_inst.gclk\[32\] dig_ctrl_inst.latch_mem_inst.RAM\[32\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_56_Right_56 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_34_56 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_1962_ VDPWR VGND VDPWR VGND net97 _0622_ dig_ctrl_inst.latch_mem_inst.RAM\[52\]\[5\]
+ net38 sky130_fd_sc_hd__and3_2
XFILLER_0_43_337 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1893_ VGND VDPWR VDPWR VGND _0525_ _0554_ _0531_ dig_ctrl_inst.latch_mem_inst.RAM\[3\]\[4\]
+ _1180_ _0526_ sky130_fd_sc_hd__a2111o_1
XPHY_EDGE_ROW_65_Right_65 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2445_ VGND VDPWR VDPWR VGND _1027_ _1022_ _1023_ _1028_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_11_267 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_2514_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.data\[5\] net151 _0040_ clknet_leaf_13_clk
+ sky130_fd_sc_hd__dfrtp_1
X_2376_ VGND VDPWR VDPWR VGND _1002_ _0996_ net339 _0065_ sky130_fd_sc_hd__mux2_1
X_1327_ VDPWR VGND VDPWR VGND _1168_ net167 net265 _1169_ sky130_fd_sc_hd__a21o_1
X_1258_ VDPWR VGND VDPWR VGND net257 _1100_ net261 dig_ctrl_inst.cpu_inst.regs\[3\]\[1\]
+ sky130_fd_sc_hd__and3_2
XPHY_EDGE_ROW_74_Right_74 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[20\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND net182 dig_ctrl_inst.latch_mem_inst.gclk\[20\] dig_ctrl_inst.latch_mem_inst.RAM\[20\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_46_153 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[58\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND net202 dig_ctrl_inst.latch_mem_inst.gclk\[58\] dig_ctrl_inst.latch_mem_inst.RAM\[58\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[61\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[61\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[61\]._gclk sky130_fd_sc_hd__clkbuf_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[47\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND net218 dig_ctrl_inst.latch_mem_inst.gclk\[47\] dig_ctrl_inst.latch_mem_inst.RAM\[47\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_20_25 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_25_337 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2230_ VGND VDPWR VDPWR VGND _0262_ _0873_ _0247_ _0841_ _0874_ sky130_fd_sc_hd__a31o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[36\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND net230 dig_ctrl_inst.latch_mem_inst.gclk\[36\] dig_ctrl_inst.latch_mem_inst.RAM\[36\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
X_2161_ VGND VDPWR VDPWR VGND _0774_ _0807_ net246 net247 sky130_fd_sc_hd__nor3_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[2\].gen_latches\[7\].p_latch VGND VDPWR VDPWR
+ VGND net179 dig_ctrl_inst.latch_mem_inst.gclk\[2\] dig_ctrl_inst.latch_mem_inst.RAM\[2\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
X_2092_ VDPWR VGND VDPWR VGND _0748_ _0711_ _0750_ _0746_ _0749_ sky130_fd_sc_hd__or4_1
X_1945_ VDPWR VGND VDPWR VGND net96 _0605_ dig_ctrl_inst.latch_mem_inst.RAM\[54\]\[5\]
+ net42 sky130_fd_sc_hd__and3_2
XFILLER_0_0_57 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_1876_ VDPWR VGND VDPWR VGND net100 _0537_ dig_ctrl_inst.latch_mem_inst.RAM\[52\]\[4\]
+ net44 sky130_fd_sc_hd__and3_2
X_2428_ VGND VDPWR VDPWR VGND _0340_ _0399_ _1016_ _0648_ _0523_ sky130_fd_sc_hd__o211ai_1
X_2359_ VDPWR VGND VDPWR VGND _0766_ _0995_ _0876_ _0879_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_34_112 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
Xdig_ctrl_inst.latch_mem_inst.gen_words\[13\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND net189 dig_ctrl_inst.latch_mem_inst.gclk\[13\] dig_ctrl_inst.latch_mem_inst.RAM\[13\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_8_Left_86 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1730_ VGND VDPWR VDPWR VGND _0394_ net122 dig_ctrl_inst.latch_mem_inst.RAM\[17\]\[1\]
+ net136 net65 sky130_fd_sc_hd__and4_1
X_1592_ VGND VDPWR VDPWR VGND net165 _0258_ net150 sky130_fd_sc_hd__nor2_1
X_1661_ VGND VDPWR VDPWR VGND _0326_ net103 dig_ctrl_inst.latch_mem_inst.RAM\[21\]\[0\]
+ net118 net62 sky130_fd_sc_hd__and4_1
X_2144_ VGND VDPWR VDPWR VGND _0790_ net140 net164 sky130_fd_sc_hd__nand2_1
X_2213_ VDPWR VGND VDPWR VGND _0793_ _0857_ _1099_ sky130_fd_sc_hd__or2_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[29\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND net238 dig_ctrl_inst.latch_mem_inst.gclk\[29\] dig_ctrl_inst.latch_mem_inst.RAM\[29\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
X_2075_ VDPWR VGND VDPWR VGND _0733_ _0124_ dig_ctrl_inst.latch_mem_inst.RAM\[13\]\[7\]
+ dig_ctrl_inst.latch_mem_inst.RAM\[19\]\[7\] _0117_ _0720_ sky130_fd_sc_hd__a221o_1
X_1859_ VDPWR VGND VDPWR VGND _0515_ _0508_ _0521_ _0513_ _0520_ sky130_fd_sc_hd__or4_1
X_1928_ VGND VDPWR VDPWR VGND _0588_ net75 dig_ctrl_inst.latch_mem_inst.RAM\[63\]\[5\]
+ net110 net44 sky130_fd_sc_hd__and4_1
XFILLER_0_8_334 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
Xdig_ctrl_inst.latch_mem_inst.gen_words\[17\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND net183 dig_ctrl_inst.latch_mem_inst.gclk\[17\] dig_ctrl_inst.latch_mem_inst.RAM\[17\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_22_104 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
Xdig_ctrl_inst.latch_mem_inst.genblk1\[39\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[39\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[39\]._gclk clknet_leaf_0_clk sky130_fd_sc_hd__dlclkp_1
XFILLER_0_26_79 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_5_337 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_5_304 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_1713_ VDPWR VGND VDPWR VGND net112 _0377_ dig_ctrl_inst.latch_mem_inst.RAM\[50\]\[1\]
+ net39 sky130_fd_sc_hd__and3_2
X_1644_ VDPWR VGND VDPWR VGND net98 _0309_ dig_ctrl_inst.latch_mem_inst.RAM\[20\]\[0\]
+ net68 sky130_fd_sc_hd__and3_2
XFILLER_0_67_42 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1575_ VGND VDPWR VDPWR VGND _0238_ _0241_ _0240_ sky130_fd_sc_hd__or2_1
X_2127_ VGND VDPWR VDPWR VGND _0773_ net247 net246 sky130_fd_sc_hd__nand2_1
X_2058_ VDPWR VGND VDPWR VGND net125 _0716_ dig_ctrl_inst.latch_mem_inst.RAM\[4\]\[7\]
+ net97 sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.genblk1\[41\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[41\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[41\]._gclk clknet_leaf_16_clk sky130_fd_sc_hd__dlclkp_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[54\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[54\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[54\]._gclk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_50_276 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_1360_ VDPWR VGND VDPWR VGND net106 _0113_ net127 net91 sky130_fd_sc_hd__and3_2
X_1291_ VDPWR VGND VDPWR VGND net257 _1133_ net261 dig_ctrl_inst.cpu_inst.regs\[3\]\[2\]
+ sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[62\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND net236 dig_ctrl_inst.latch_mem_inst.gclk\[62\] dig_ctrl_inst.latch_mem_inst.RAM\[62\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
X_1489_ VDPWR VGND VDPWR VGND dig_ctrl_inst.spi_receiver_inst.spi_cnt\[0\] dig_ctrl_inst.spi_receiver_inst.spi_cnt\[1\]
+ _0179_ _0177_ sky130_fd_sc_hd__a21oi_1
X_1627_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[10\]\[0\] _1190_ _0292_
+ dig_ctrl_inst.latch_mem_inst.RAM\[31\]\[0\] _0133_ sky130_fd_sc_hd__a22o_1
X_1558_ VGND VDPWR VDPWR VGND _0224_ _0222_ _0223_ sky130_fd_sc_hd__and2b_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[50\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND net179 dig_ctrl_inst.latch_mem_inst.gclk\[50\] dig_ctrl_inst.latch_mem_inst.RAM\[50\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_2_3 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_21_Left_99 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2530_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[1\]\[2\] net153 _0056_
+ clknet_leaf_11_clk sky130_fd_sc_hd__dfrtp_1
X_2392_ VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_receiver_inst.spi_cnt\[0\] dig_ctrl_inst.spi_data_i\[2\]
+ dig_ctrl_inst.spi_data_i\[3\] _1006_ sky130_fd_sc_hd__mux2_1
X_2461_ VGND VDPWR VDPWR VGND dig_ctrl_inst.synchronizer_port_i_inst\[7\].out net169
+ net296 clknet_leaf_4_clk sky130_fd_sc_hd__dfrtp_1
X_1343_ VGND VDPWR VDPWR VGND _1139_ _1181_ _1122_ sky130_fd_sc_hd__nor2_1
X_1412_ VDPWR VGND VDPWR VGND net98 dig_ctrl_inst.latch_mem_inst.data_we\[36\] net147
+ net56 sky130_fd_sc_hd__and3_2
Xwire36 VGND VDPWR VDPWR VGND net36 _0690_ sky130_fd_sc_hd__clkbuf_1
X_1274_ VDPWR VGND VDPWR VGND net257 _1116_ net261 dig_ctrl_inst.cpu_inst.regs\[3\]\[3\]
+ sky130_fd_sc_hd__and3_2
XFILLER_0_3_57 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_16_clk VGND VDPWR VDPWR VGND clknet_leaf_16_clk clknet_1_0__leaf_clk
+ sky130_fd_sc_hd__clkbuf_8
Xfanout167 VDPWR VGND VDPWR VGND net167 _1082_ sky130_fd_sc_hd__buf_2
Xfanout156 VGND VDPWR VDPWR VGND net156 net157 sky130_fd_sc_hd__clkbuf_4
Xfanout101 VDPWR VGND VDPWR VGND net101 net102 sky130_fd_sc_hd__buf_2
Xfanout145 VGND VDPWR VDPWR VGND net146 net145 sky130_fd_sc_hd__clkbuf_2
Xfanout189 VDPWR VGND VDPWR VGND net189 net284 sky130_fd_sc_hd__buf_2
Xfanout178 VGND VDPWR VDPWR VGND net185 net178 sky130_fd_sc_hd__clkbuf_2
Xfanout112 VGND VDPWR VDPWR VGND net113 net112 sky130_fd_sc_hd__clkbuf_2
Xfanout134 VGND VDPWR VDPWR VGND net135 net134 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_64_187 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[43\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND net186 dig_ctrl_inst.latch_mem_inst.gclk\[43\] dig_ctrl_inst.latch_mem_inst.RAM\[43\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_34_46 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1892_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[17\]\[4\] _0122_ _0553_
+ dig_ctrl_inst.latch_mem_inst.RAM\[42\]\[4\] _0145_ sky130_fd_sc_hd__a22o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[32\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND net205 dig_ctrl_inst.latch_mem_inst.gclk\[32\] dig_ctrl_inst.latch_mem_inst.RAM\[32\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
X_1961_ VGND VDPWR VDPWR VGND _0621_ net104 dig_ctrl_inst.latch_mem_inst.RAM\[35\]\[5\]
+ net138 net48 sky130_fd_sc_hd__and4_1
XFILLER_0_50_89 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
X_2513_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.data\[4\] net151 _0039_ clknet_leaf_14_clk
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_5_clk VGND VDPWR VDPWR VGND clknet_leaf_5_clk clknet_1_1__leaf_clk sky130_fd_sc_hd__clkbuf_8
X_2444_ VDPWR VGND VDPWR VGND dig_ctrl_inst.spi_addr\[1\] _1027_ dig_ctrl_inst.spi_addr\[0\]
+ dig_ctrl_inst.spi_addr\[2\] sky130_fd_sc_hd__and3_2
X_1326_ VGND VDPWR VDPWR VGND _1061_ _1164_ _1165_ _1166_ _1167_ _1168_ sky130_fd_sc_hd__o41a_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[21\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND net222 dig_ctrl_inst.latch_mem_inst.gclk\[21\] dig_ctrl_inst.latch_mem_inst.RAM\[21\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
X_2375_ VGND VDPWR VDPWR VGND _1002_ _0995_ net320 _0064_ sky130_fd_sc_hd__mux2_1
X_1257_ VGND VDPWR VDPWR VGND _1099_ _1097_ _1096_ sky130_fd_sc_hd__nand2_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[47\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[47\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[47\]._gclk sky130_fd_sc_hd__clkbuf_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[59\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND net242 dig_ctrl_inst.latch_mem_inst.gclk\[59\] dig_ctrl_inst.latch_mem_inst.RAM\[59\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[10\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND net236 dig_ctrl_inst.latch_mem_inst.gclk\[10\] dig_ctrl_inst.latch_mem_inst.RAM\[10\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[47\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND net182 dig_ctrl_inst.latch_mem_inst.gclk\[47\] dig_ctrl_inst.latch_mem_inst.RAM\[47\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[3\].gen_latches\[2\].p_latch VGND VDPWR VDPWR
+ VGND net222 dig_ctrl_inst.latch_mem_inst.gclk\[3\] dig_ctrl_inst.latch_mem_inst.RAM\[3\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_29_57 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_2160_ VGND VDPWR VDPWR VGND _1039_ net247 _0804_ _0806_ sky130_fd_sc_hd__or3b_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[36\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND net197 dig_ctrl_inst.latch_mem_inst.gclk\[36\] dig_ctrl_inst.latch_mem_inst.RAM\[36\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
X_2091_ VGND VDPWR VDPWR VGND _0715_ _0749_ _0719_ dig_ctrl_inst.latch_mem_inst.RAM\[25\]\[7\]
+ _0129_ _0716_ sky130_fd_sc_hd__a2111o_1
X_1944_ VGND VDPWR VDPWR VGND _0604_ net129 dig_ctrl_inst.latch_mem_inst.RAM\[3\]\[5\]
+ net137 net108 sky130_fd_sc_hd__and4_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[25\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND net212 dig_ctrl_inst.latch_mem_inst.gclk\[25\] dig_ctrl_inst.latch_mem_inst.RAM\[25\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_9_23 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_1875_ VDPWR VGND VDPWR VGND net125 _0536_ dig_ctrl_inst.latch_mem_inst.RAM\[6\]\[4\]
+ net93 sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_input_latches\[3\].n_latch VGND VDPWR VDPWR VGND
+ dig_ctrl_inst.data_out\[3\] clknet_leaf_9_clk dig_ctrl_inst.latch_mem_inst.wdata\[3\]
+ sky130_fd_sc_hd__dlxtn_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[46\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[46\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[46\]._gclk clknet_leaf_18_clk sky130_fd_sc_hd__dlclkp_1
XFILLER_0_3_221 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2427_ VGND VDPWR VDPWR VGND _1015_ _1014_ _0195_ sky130_fd_sc_hd__nand2_1
X_1309_ VDPWR VGND VDPWR VGND net262 _1151_ net259 dig_ctrl_inst.cpu_inst.regs\[0\]\[5\]
+ sky130_fd_sc_hd__or3_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[14\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND net234 dig_ctrl_inst.latch_mem_inst.gclk\[14\] dig_ctrl_inst.latch_mem_inst.RAM\[14\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_19_90 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_2289_ VGND VDPWR VDPWR VGND _0930_ net159 _1147_ sky130_fd_sc_hd__nand2_1
X_2358_ VGND VDPWR VDPWR VGND _0991_ _0994_ net332 _0055_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_198 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
Xdig_ctrl_inst.latch_mem_inst.gen_words\[7\].gen_latches\[3\].p_latch VGND VDPWR VDPWR
+ VGND net218 dig_ctrl_inst.latch_mem_inst.gclk\[7\] dig_ctrl_inst.latch_mem_inst.RAM\[7\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_25_113 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1660_ VGND VDPWR VDPWR VGND _0322_ _0325_ _0324_ dig_ctrl_inst.latch_mem_inst.RAM\[57\]\[0\]
+ _0157_ _0323_ sky130_fd_sc_hd__a2111o_1
Xwire162 VGND VDPWR VDPWR VGND _1130_ net162 sky130_fd_sc_hd__clkbuf_2
X_1591_ VGND VDPWR VDPWR VGND _0257_ _0247_ _0241_ sky130_fd_sc_hd__nand2_1
X_2143_ VGND VDPWR VDPWR VGND _0788_ _0789_ net150 sky130_fd_sc_hd__nor2_1
X_2212_ VGND VDPWR VDPWR VGND _0771_ dig_ctrl_inst.cpu_inst.regs\[0\]\[1\] _0856_
+ _0047_ sky130_fd_sc_hd__mux2_1
X_2074_ VDPWR VGND VDPWR VGND _0732_ _0159_ dig_ctrl_inst.latch_mem_inst.RAM\[22\]\[7\]
+ dig_ctrl_inst.latch_mem_inst.RAM\[59\]\[7\] _0127_ _0731_ sky130_fd_sc_hd__a221o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[29\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND net206 dig_ctrl_inst.latch_mem_inst.gclk\[29\] dig_ctrl_inst.latch_mem_inst.RAM\[29\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_31_149 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_1858_ VDPWR VGND VDPWR VGND _0518_ _0516_ _0520_ _0517_ _0519_ sky130_fd_sc_hd__or4_1
X_1927_ VGND VDPWR VDPWR VGND _0587_ net89 dig_ctrl_inst.latch_mem_inst.RAM\[57\]\[5\]
+ net117 net37 sky130_fd_sc_hd__and4_1
X_1789_ VDPWR VGND VDPWR VGND net82 _0452_ dig_ctrl_inst.latch_mem_inst.RAM\[26\]\[2\]
+ net66 sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[18\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND net219 dig_ctrl_inst.latch_mem_inst.gclk\[18\] dig_ctrl_inst.latch_mem_inst.RAM\[18\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
X_2609__273 VGND VDPWR VDPWR VGND net273 _2609__273/HI sky130_fd_sc_hd__conb_1
XFILLER_0_30_160 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
Xhold70 VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[1\]\[0\] net352 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_1 VGND VDPWR VDPWR VGND _0098_ sky130_fd_sc_hd__diode_2
X_1643_ VDPWR VGND VDPWR VGND net82 _0308_ dig_ctrl_inst.latch_mem_inst.RAM\[42\]\[0\]
+ net57 sky130_fd_sc_hd__and3_2
X_1712_ VDPWR VGND VDPWR VGND net84 _0376_ dig_ctrl_inst.latch_mem_inst.RAM\[24\]\[1\]
+ net59 sky130_fd_sc_hd__and3_2
XFILLER_0_13_127 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1574_ VGND VDPWR VDPWR VGND net163 _0240_ _1113_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_46 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2057_ VDPWR VGND VDPWR VGND net112 _0715_ dig_ctrl_inst.latch_mem_inst.RAM\[50\]\[7\]
+ net40 sky130_fd_sc_hd__and3_2
X_2126_ VDPWR VGND VDPWR VGND _0189_ _0770_ _0768_ net177 _0772_ sky130_fd_sc_hd__o211a_2
XFILLER_0_44_263 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1290_ VDPWR VGND VDPWR VGND net261 _1132_ net257 dig_ctrl_inst.cpu_inst.regs\[0\]\[2\]
+ sky130_fd_sc_hd__or3_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[62\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND net205 dig_ctrl_inst.latch_mem_inst.gclk\[62\] dig_ctrl_inst.latch_mem_inst.RAM\[62\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
X_1626_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[27\]\[0\] _0130_ _0291_
+ dig_ctrl_inst.latch_mem_inst.RAM\[60\]\[0\] _0160_ sky130_fd_sc_hd__a22o_1
X_1488_ VDPWR VGND VDPWR VGND dig_ctrl_inst.spi_receiver_inst.spi_cnt\[1\] _0178_
+ dig_ctrl_inst.spi_receiver_inst.spi_cnt\[0\] _0177_ sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[51\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND net224 dig_ctrl_inst.latch_mem_inst.gclk\[51\] dig_ctrl_inst.latch_mem_inst.RAM\[51\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
X_1557_ VGND VDPWR VDPWR VGND _0223_ _0221_ _0172_ sky130_fd_sc_hd__nand2_1
X_2109_ VGND VDPWR VDPWR VGND _0762_ _0522_ dig_ctrl_inst.cpu_inst.data\[3\] _0038_
+ sky130_fd_sc_hd__mux2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[40\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND net236 dig_ctrl_inst.latch_mem_inst.gclk\[40\] dig_ctrl_inst.latch_mem_inst.RAM\[40\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
X_2460_ VGND VDPWR VDPWR VGND dig_ctrl_inst.synchronizer_port_i_inst\[7\].pipe\[0\]
+ net168 net10 clknet_leaf_4_clk sky130_fd_sc_hd__dfrtp_1
X_2391_ VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_receiver_inst.spi_cnt\[0\] dig_ctrl_inst.spi_data_i\[6\]
+ _1005_ dig_ctrl_inst.spi_receiver_inst.spi_cnt\[1\] dig_ctrl_inst.spi_data_i\[5\]
+ dig_ctrl_inst.spi_data_i\[7\] dig_ctrl_inst.spi_data_i\[4\] sky130_fd_sc_hd__mux4_1
X_1342_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[3\] _1180_ net146
+ sky130_fd_sc_hd__and2_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[11\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[11\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[11\]._gclk sky130_fd_sc_hd__clkbuf_4
X_1411_ VDPWR VGND VDPWR VGND _0139_ net52 _1182_ sky130_fd_sc_hd__and2_1
X_1273_ VGND VDPWR VDPWR VGND _1056_ _1071_ _1115_ _1114_ sky130_fd_sc_hd__or3_2
XFILLER_0_58_141 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_174 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
Xfanout113 VGND VDPWR VDPWR VGND net113 _1177_ sky130_fd_sc_hd__clkbuf_4
X_2589_ VGND VDPWR VDPWR VGND net23 net174 _0103_ clknet_leaf_6_clk sky130_fd_sc_hd__dfrtp_1
Xfanout102 VGND VDPWR VDPWR VGND net102 net103 sky130_fd_sc_hd__clkbuf_4
X_1609_ VDPWR VGND VDPWR VGND _0135_ _0127_ _0274_ _0128_ _0136_ sky130_fd_sc_hd__or4_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[55\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND net213 dig_ctrl_inst.latch_mem_inst.gclk\[55\] dig_ctrl_inst.latch_mem_inst.RAM\[55\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_14_299 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xfanout168 VGND VDPWR VDPWR VGND net168 net170 sky130_fd_sc_hd__clkbuf_4
Xfanout135 VDPWR VGND VDPWR VGND net135 _1141_ sky130_fd_sc_hd__buf_2
Xfanout157 VGND VDPWR VDPWR VGND net157 dig_ctrl_inst.cpu_inst.rst_ni sky130_fd_sc_hd__clkbuf_4
Xfanout146 VGND VDPWR VDPWR VGND net148 net146 sky130_fd_sc_hd__clkbuf_2
Xfanout124 VGND VDPWR VDPWR VGND net126 net124 sky130_fd_sc_hd__clkbuf_2
Xfanout179 VGND VDPWR VDPWR VGND net180 net179 sky130_fd_sc_hd__clkbuf_2
Xdig_ctrl_inst.latch_mem_inst.genblk1\[53\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[53\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[53\]._gclk clknet_leaf_19_clk sky130_fd_sc_hd__dlclkp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[44\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND net228 dig_ctrl_inst.latch_mem_inst.gclk\[44\] dig_ctrl_inst.latch_mem_inst.RAM\[44\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_9_271 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_1960_ VGND VDPWR VDPWR VGND _0620_ net79 dig_ctrl_inst.latch_mem_inst.RAM\[45\]\[5\]
+ net120 net55 sky130_fd_sc_hd__and4_1
X_1891_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[1\]\[4\] _1175_ _0552_
+ dig_ctrl_inst.latch_mem_inst.RAM\[57\]\[4\] _0157_ sky130_fd_sc_hd__a22o_1
X_2443_ VDPWR VGND VDPWR VGND _1026_ _1042_ _1023_ _1024_ _0108_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_11_225 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_2512_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.data\[3\] net151 _0038_ clknet_leaf_10_clk
+ sky130_fd_sc_hd__dfrtp_1
X_1325_ VDPWR VGND VDPWR VGND net262 _1167_ net258 dig_ctrl_inst.cpu_inst.regs\[0\]\[4\]
+ sky130_fd_sc_hd__or3_1
X_1256_ VGND VDPWR VDPWR VGND _1063_ _1093_ _1094_ _1095_ _1097_ _1098_ sky130_fd_sc_hd__o41a_4
X_2374_ VGND VDPWR VDPWR VGND _1002_ _0994_ net325 _0063_ sky130_fd_sc_hd__mux2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[21\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND net186 dig_ctrl_inst.latch_mem_inst.gclk\[21\] dig_ctrl_inst.latch_mem_inst.RAM\[21\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_49_Left_127 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[59\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND net210 dig_ctrl_inst.latch_mem_inst.gclk\[59\] dig_ctrl_inst.latch_mem_inst.RAM\[59\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[10\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND net203 dig_ctrl_inst.latch_mem_inst.gclk\[10\] dig_ctrl_inst.latch_mem_inst.RAM\[10\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_58_Left_136 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[48\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND net221 dig_ctrl_inst.latch_mem_inst.gclk\[48\] dig_ctrl_inst.latch_mem_inst.RAM\[48\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_67_Left_145 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_76_Left_154 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[37\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND net238 dig_ctrl_inst.latch_mem_inst.gclk\[37\] dig_ctrl_inst.latch_mem_inst.RAM\[37\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[3\].gen_latches\[6\].p_latch VGND VDPWR VDPWR
+ VGND net189 dig_ctrl_inst.latch_mem_inst.gclk\[3\] dig_ctrl_inst.latch_mem_inst.RAM\[3\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
X_2090_ VGND VDPWR VDPWR VGND _0712_ _0748_ _0730_ dig_ctrl_inst.latch_mem_inst.RAM\[35\]\[7\]
+ _0138_ _0714_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_45_57 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_0_15 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_1943_ VGND VDPWR VDPWR VGND _0603_ net78 dig_ctrl_inst.latch_mem_inst.RAM\[29\]\[5\]
+ net121 net68 sky130_fd_sc_hd__and4_1
X_1874_ VDPWR VGND VDPWR VGND net100 _0535_ dig_ctrl_inst.latch_mem_inst.RAM\[36\]\[4\]
+ net54 sky130_fd_sc_hd__and3_2
XFILLER_0_43_147 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_9_35 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_2426_ VGND VDPWR VDPWR VGND _1014_ dig_ctrl_inst.stb_dd dig_ctrl_inst.cpu_inst.cpu_state\[2\]
+ net167 sky130_fd_sc_hd__a21bo_1
Xdig_ctrl_inst.latch_mem_inst.gen_input_latches\[7\].n_latch VGND VDPWR VDPWR VGND
+ dig_ctrl_inst.data_out\[7\] clknet_leaf_9_clk dig_ctrl_inst.latch_mem_inst.wdata\[7\]
+ sky130_fd_sc_hd__dlxtn_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[25\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND net180 dig_ctrl_inst.latch_mem_inst.gclk\[25\] dig_ctrl_inst.latch_mem_inst.RAM\[25\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
X_1308_ VGND VDPWR VDPWR VGND _1150_ net259 dig_ctrl_inst.cpu_inst.regs\[1\]\[5\]
+ sky130_fd_sc_hd__and2b_1
X_1239_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[0\]\[0\] _1081_ net176
+ _1078_ _1079_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_36_3 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_2288_ VGND VDPWR VDPWR VGND _1147_ _0929_ net159 sky130_fd_sc_hd__or2_1
X_2357_ VDPWR VGND VDPWR VGND _0853_ _0839_ _0994_ _0842_ _0993_ sky130_fd_sc_hd__or4_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[14\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND net199 dig_ctrl_inst.latch_mem_inst.gclk\[14\] dig_ctrl_inst.latch_mem_inst.RAM\[14\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[7\].gen_latches\[7\].p_latch VGND VDPWR VDPWR
+ VGND net184 dig_ctrl_inst.latch_mem_inst.gclk\[7\] dig_ctrl_inst.latch_mem_inst.RAM\[7\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_0_225 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_1590_ VGND VDPWR VDPWR VGND _0254_ _1039_ _0253_ _0255_ _0256_ sky130_fd_sc_hd__a31o_1
X_2073_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[37\]\[7\] _0140_ _0731_
+ dig_ctrl_inst.latch_mem_inst.RAM\[39\]\[7\] _0142_ sky130_fd_sc_hd__a22o_1
X_2142_ VGND VDPWR VDPWR VGND _0788_ net140 net165 sky130_fd_sc_hd__nand2_1
X_2211_ VDPWR VGND VDPWR VGND _0853_ _0839_ _0856_ _0842_ _0855_ sky130_fd_sc_hd__or4_1
X_1788_ VGND VDPWR VDPWR VGND _0448_ _0451_ _0450_ dig_ctrl_inst.latch_mem_inst.RAM\[35\]\[2\]
+ _0138_ _0449_ sky130_fd_sc_hd__a2111o_1
X_1857_ VGND VDPWR VDPWR VGND _0467_ _0519_ _0490_ dig_ctrl_inst.latch_mem_inst.RAM\[5\]\[3\]
+ _0272_ _0480_ sky130_fd_sc_hd__a2111o_1
X_1926_ VDPWR VGND VDPWR VGND net133 _0586_ dig_ctrl_inst.latch_mem_inst.RAM\[48\]\[5\]
+ net37 sky130_fd_sc_hd__and3_2
X_2409_ VGND VDPWR VDPWR VGND _1012_ dig_ctrl_inst.cpu_inst.port_o\[0\] net25 _0088_
+ sky130_fd_sc_hd__mux2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[18\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND net192 dig_ctrl_inst.latch_mem_inst.gclk\[18\] dig_ctrl_inst.latch_mem_inst.RAM\[18\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
Xhold60 VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[3\]\[0\] net342 sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[3\]\[3\] net353 sky130_fd_sc_hd__dlygate4sd3_1
X_1642_ VDPWR VGND VDPWR VGND net113 _0307_ dig_ctrl_inst.latch_mem_inst.RAM\[50\]\[0\]
+ net46 sky130_fd_sc_hd__and3_2
XANTENNA_2 VGND VDPWR VDPWR VGND _0115_ sky130_fd_sc_hd__diode_2
X_1711_ VDPWR VGND VDPWR VGND _0375_ _0152_ dig_ctrl_inst.latch_mem_inst.RAM\[45\]\[1\]
+ dig_ctrl_inst.latch_mem_inst.RAM\[49\]\[1\] _0147_ _0374_ sky130_fd_sc_hd__a221o_1
X_1573_ VGND VDPWR VDPWR VGND _0239_ net163 _1113_ sky130_fd_sc_hd__nand2_1
X_2056_ VDPWR VGND VDPWR VGND net134 _0714_ dig_ctrl_inst.latch_mem_inst.RAM\[32\]\[7\]
+ net50 sky130_fd_sc_hd__and3_2
X_2125_ VGND VDPWR VDPWR VGND net177 _0770_ _0768_ _0189_ _0771_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_44_253 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1909_ VGND VDPWR VDPWR VGND _0538_ _0570_ _0541_ dig_ctrl_inst.latch_mem_inst.RAM\[35\]\[4\]
+ _0138_ _0540_ sky130_fd_sc_hd__a2111o_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[58\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[58\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[58\]._gclk clknet_leaf_16_clk sky130_fd_sc_hd__dlclkp_1
XFILLER_0_50_212 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_35_264 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
Xdig_ctrl_inst.latch_mem_inst.genblk1\[60\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[60\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[60\]._gclk clknet_leaf_17_clk sky130_fd_sc_hd__dlclkp_1
XFILLER_0_53_57 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1625_ VGND VDPWR VDPWR VGND _0287_ _0290_ _0289_ dig_ctrl_inst.latch_mem_inst.RAM\[3\]\[0\]
+ _1180_ _0288_ sky130_fd_sc_hd__a2111o_1
X_1556_ VGND VDPWR VDPWR VGND _0221_ _0222_ _0172_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_320 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_1487_ VGND VDPWR VDPWR VGND _0176_ _0001_ dig_ctrl_inst.spi_receiver_inst.spi_cnt\[0\]
+ sky130_fd_sc_hd__xnor2_1
X_2039_ VGND VDPWR VDPWR VGND _0695_ _0698_ _0697_ dig_ctrl_inst.latch_mem_inst.RAM\[7\]\[6\]
+ _1184_ _0696_ sky130_fd_sc_hd__a2111o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[51\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND net190 dig_ctrl_inst.latch_mem_inst.gclk\[51\] dig_ctrl_inst.latch_mem_inst.RAM\[51\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_30_Left_108 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2108_ VGND VDPWR VDPWR VGND _0762_ _0462_ dig_ctrl_inst.cpu_inst.data\[2\] _0037_
+ sky130_fd_sc_hd__mux2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[40\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND net203 dig_ctrl_inst.latch_mem_inst.gclk\[40\] dig_ctrl_inst.latch_mem_inst.RAM\[40\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_4_191 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.genblk1\[50\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[50\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[50\]._gclk sky130_fd_sc_hd__clkbuf_4
X_1410_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[35\] _0138_ net143
+ sky130_fd_sc_hd__and2_1
X_2390_ VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_receiver_inst.spi_cs_sync dig_ctrl_inst.spi_receiver_inst.spi_sclk_sync
+ _1004_ dig_ctrl_inst.spi_receiver_inst.spi_sclk_delayed sky130_fd_sc_hd__or3b_1
X_1341_ VGND VDPWR VDPWR VGND net136 net130 net109 _1180_ sky130_fd_sc_hd__and3_4
X_1272_ VGND VDPWR VDPWR VGND _1114_ _1111_ _1110_ _1109_ net176 _1112_ sky130_fd_sc_hd__a41o_4
XFILLER_0_58_153 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xfanout147 VGND VDPWR VDPWR VGND net148 net147 sky130_fd_sc_hd__clkbuf_2
X_2588_ VGND VDPWR VDPWR VGND net22 net174 _0102_ clknet_leaf_6_clk sky130_fd_sc_hd__dfrtp_1
Xfanout136 VGND VDPWR VDPWR VGND net136 _1140_ sky130_fd_sc_hd__clkbuf_4
Xfanout103 VGND VDPWR VDPWR VGND net103 _1181_ sky130_fd_sc_hd__clkbuf_4
Xfanout114 VDPWR VGND VDPWR VGND net114 _1176_ sky130_fd_sc_hd__buf_2
X_1608_ VDPWR VGND VDPWR VGND _0119_ _1178_ _0273_ _1187_ _0272_ sky130_fd_sc_hd__or4_1
X_1539_ VDPWR VGND VDPWR VGND dig_ctrl_inst.cpu_inst.ip\[2\] _0205_ _0022_ _0197_
+ _0208_ sky130_fd_sc_hd__a22o_1
Xfanout125 VDPWR VGND VDPWR VGND net125 net126 sky130_fd_sc_hd__buf_2
Xfanout169 VGND VDPWR VDPWR VGND net169 net170 sky130_fd_sc_hd__clkbuf_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[55\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND net181 dig_ctrl_inst.latch_mem_inst.gclk\[55\] dig_ctrl_inst.latch_mem_inst.RAM\[55\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
Xfanout158 VDPWR VGND VDPWR VGND net158 _1168_ sky130_fd_sc_hd__buf_2
XFILLER_0_64_112 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[44\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND net197 dig_ctrl_inst.latch_mem_inst.gclk\[44\] dig_ctrl_inst.latch_mem_inst.RAM\[44\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[0\].gen_latches\[0\].p_latch VGND VDPWR VDPWR
+ VGND net239 dig_ctrl_inst.latch_mem_inst.gclk\[0\] dig_ctrl_inst.latch_mem_inst.RAM\[0\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[33\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND net217 dig_ctrl_inst.latch_mem_inst.gclk\[33\] dig_ctrl_inst.latch_mem_inst.RAM\[33\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_16_Right_16 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[22\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND net233 dig_ctrl_inst.latch_mem_inst.gclk\[22\] dig_ctrl_inst.latch_mem_inst.RAM\[22\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
X_1890_ VGND VDPWR VDPWR VGND _0524_ _0551_ _0533_ dig_ctrl_inst.latch_mem_inst.RAM\[55\]\[4\]
+ _0155_ _0532_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_70_137 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_25_Right_25 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2442_ VDPWR VGND VDPWR VGND dig_ctrl_inst.spi_addr\[1\] dig_ctrl_inst.spi_addr\[0\]
+ _1022_ _1026_ sky130_fd_sc_hd__a21o_1
X_2373_ VGND VDPWR VDPWR VGND _1002_ _0992_ net326 _0062_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_11 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_11_237 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_2511_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.data\[2\] net152 _0037_ clknet_leaf_10_clk
+ sky130_fd_sc_hd__dfrtp_1
X_1324_ VGND VDPWR VDPWR VGND _1166_ net258 dig_ctrl_inst.cpu_inst.regs\[1\]\[4\]
+ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_34_Right_34 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1255_ VDPWR VGND VDPWR VGND net253 _1097_ net249 dig_ctrl_inst.cpu_inst.regs\[0\]\[1\]
+ sky130_fd_sc_hd__or3_1
XFILLER_0_19_337 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_43_Right_43 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_6_253 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_52_Right_52 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2603__269 VGND VDPWR VDPWR VGND net269 _2603__269/HI sky130_fd_sc_hd__conb_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[4\].gen_latches\[1\].p_latch VGND VDPWR VDPWR
+ VGND net235 dig_ctrl_inst.latch_mem_inst.gclk\[4\] dig_ctrl_inst.latch_mem_inst.RAM\[4\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_4_91 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[48\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND net186 dig_ctrl_inst.latch_mem_inst.gclk\[48\] dig_ctrl_inst.latch_mem_inst.RAM\[48\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_61_Right_61 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_20_17 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_70_Right_70 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[37\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND net207 dig_ctrl_inst.latch_mem_inst.gclk\[37\] dig_ctrl_inst.latch_mem_inst.RAM\[37\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_45_25 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
Xdig_ctrl_inst.latch_mem_inst.gen_words\[26\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND net224 dig_ctrl_inst.latch_mem_inst.gclk\[26\] dig_ctrl_inst.latch_mem_inst.RAM\[26\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_28_156 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1942_ VDPWR VGND VDPWR VGND net97 _0602_ dig_ctrl_inst.latch_mem_inst.RAM\[36\]\[5\]
+ net49 sky130_fd_sc_hd__and3_2
XFILLER_0_51_181 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_1873_ VDPWR VGND VDPWR VGND net134 _0534_ dig_ctrl_inst.latch_mem_inst.RAM\[32\]\[4\]
+ net50 sky130_fd_sc_hd__and3_2
X_2425_ VGND VDPWR VDPWR VGND _1013_ dig_ctrl_inst.cpu_inst.port_o\[7\] net311 _0103_
+ sky130_fd_sc_hd__mux2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[15\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND net241 dig_ctrl_inst.latch_mem_inst.gclk\[15\] dig_ctrl_inst.latch_mem_inst.RAM\[15\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
X_2356_ VGND VDPWR VDPWR VGND _0851_ _0993_ _0766_ sky130_fd_sc_hd__nor2_1
X_2287_ VDPWR VGND VDPWR VGND _0050_ _0928_ _0771_ _0923_ _0772_ net341 sky130_fd_sc_hd__o32a_1
X_1307_ VDPWR VGND VDPWR VGND net259 _1149_ net263 dig_ctrl_inst.cpu_inst.regs\[3\]\[5\]
+ sky130_fd_sc_hd__and3_2
X_1238_ VGND VDPWR VDPWR VGND net176 _1080_ _1078_ dig_ctrl_inst.cpu_inst.regs\[0\]\[0\]
+ _1079_ sky130_fd_sc_hd__o22a_2
XFILLER_0_29_3 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_34_137 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[8\].gen_latches\[2\].p_latch VGND VDPWR VDPWR
+ VGND net224 dig_ctrl_inst.latch_mem_inst.gclk\[8\] dig_ctrl_inst.latch_mem_inst.RAM\[8\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[43\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[43\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[43\]._gclk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_15_17 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_0_237 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
X_2210_ VGND VDPWR VDPWR VGND _0854_ _0767_ _0851_ _0855_ _0768_ sky130_fd_sc_hd__a2bb2o_1
X_2141_ VGND VDPWR VDPWR VGND _0781_ _0787_ _0782_ _0776_ _0786_ sky130_fd_sc_hd__o22a_1
X_2072_ VDPWR VGND VDPWR VGND net125 _0730_ dig_ctrl_inst.latch_mem_inst.RAM\[2\]\[7\]
+ net112 sky130_fd_sc_hd__and3_2
X_1925_ VDPWR VGND VDPWR VGND net124 _0585_ dig_ctrl_inst.latch_mem_inst.RAM\[8\]\[5\]
+ net84 sky130_fd_sc_hd__and3_2
XFILLER_0_16_137 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1787_ VDPWR VGND VDPWR VGND net87 _0450_ dig_ctrl_inst.latch_mem_inst.RAM\[56\]\[2\]
+ net45 sky130_fd_sc_hd__and3_2
X_1856_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[19\]\[3\] _0124_ _0518_
+ dig_ctrl_inst.latch_mem_inst.RAM\[57\]\[3\] _0157_ sky130_fd_sc_hd__a22o_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[19\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND net231 dig_ctrl_inst.latch_mem_inst.gclk\[19\] dig_ctrl_inst.latch_mem_inst.RAM\[19\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
X_2408_ VDPWR VGND VDPWR VGND _1012_ _0824_ _0187_ sky130_fd_sc_hd__and2b_2
X_2339_ VGND VDPWR VDPWR VGND _0810_ _0978_ _0223_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_2_Right_2 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xhold61 VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[0\]\[5\] net343 sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[0\]\[6\] net354 sky130_fd_sc_hd__dlygate4sd3_1
Xhold50 VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[1\]\[1\] net332 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_284 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_1710_ VDPWR VGND VDPWR VGND net127 _0374_ dig_ctrl_inst.latch_mem_inst.RAM\[12\]\[1\]
+ net73 sky130_fd_sc_hd__and3_2
XANTENNA_3 VGND VDPWR VDPWR VGND _0128_ sky130_fd_sc_hd__diode_2
X_1641_ VGND VDPWR VDPWR VGND _0305_ _0298_ _0306_ _0286_ _0293_ sky130_fd_sc_hd__nor4_1
X_1572_ VDPWR VGND VDPWR VGND _0238_ net163 _1113_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_15 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
X_2124_ VDPWR VGND VDPWR VGND _1069_ _1065_ _0769_ _0770_ sky130_fd_sc_hd__a21o_1
X_2055_ VGND VDPWR VDPWR VGND _0713_ net119 dig_ctrl_inst.latch_mem_inst.RAM\[49\]\[7\]
+ net136 net43 sky130_fd_sc_hd__and4_1
X_1908_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[18\]\[4\] _0123_ _0569_
+ dig_ctrl_inst.latch_mem_inst.RAM\[45\]\[4\] _0147_ sky130_fd_sc_hd__a22o_1
X_1839_ VGND VDPWR VDPWR VGND _0477_ _0501_ _0484_ dig_ctrl_inst.latch_mem_inst.RAM\[55\]\[3\]
+ _0155_ _0482_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_35_221 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_35_276 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[63\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND net212 dig_ctrl_inst.latch_mem_inst.gclk\[63\] dig_ctrl_inst.latch_mem_inst.RAM\[63\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[52\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND net233 dig_ctrl_inst.latch_mem_inst.gclk\[52\] dig_ctrl_inst.latch_mem_inst.RAM\[52\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
X_1555_ VGND VDPWR VDPWR VGND _0221_ _0220_ net262 net258 dig_ctrl_inst.cpu_inst.regs\[0\]\[7\]
+ _0219_ sky130_fd_sc_hd__o32a_4
X_1624_ VGND VDPWR VDPWR VGND _0289_ net101 dig_ctrl_inst.latch_mem_inst.RAM\[39\]\[0\]
+ net109 net55 sky130_fd_sc_hd__and4_1
XFILLER_0_1_332 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1486_ VDPWR VGND VDPWR VGND _0176_ _0177_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_19_clk VGND VDPWR VDPWR VGND clknet_leaf_19_clk clknet_1_1__leaf_clk
+ sky130_fd_sc_hd__clkbuf_8
X_2107_ VGND VDPWR VDPWR VGND _0762_ _0399_ dig_ctrl_inst.cpu_inst.data\[1\] _0036_
+ sky130_fd_sc_hd__mux2_1
X_2038_ VGND VDPWR VDPWR VGND _0697_ net121 dig_ctrl_inst.latch_mem_inst.RAM\[33\]\[6\]
+ net137 net56 sky130_fd_sc_hd__and4_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[36\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[36\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[36\]._gclk sky130_fd_sc_hd__clkbuf_4
X_1340_ VGND VDPWR VDPWR VGND _1107_ _1179_ _1052_ _1090_ sky130_fd_sc_hd__nor3_1
X_1271_ VGND VDPWR VDPWR VGND _1112_ _1109_ net176 _1111_ _1110_ _1113_ sky130_fd_sc_hd__a41oi_4
XFILLER_0_58_165 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_73_113 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_8_clk VGND VDPWR VDPWR VGND clknet_leaf_8_clk clknet_1_1__leaf_clk sky130_fd_sc_hd__clkbuf_8
Xdig_ctrl_inst.latch_mem_inst.gen_words\[56\].gen_latches\[2\].p_latch VGND VDPWR
+ VDPWR VGND net225 dig_ctrl_inst.latch_mem_inst.gclk\[56\] dig_ctrl_inst.latch_mem_inst.RAM\[56\]\[2\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_14_257 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xfanout104 VDPWR VGND VDPWR VGND net104 net105 sky130_fd_sc_hd__buf_2
Xfanout126 VGND VDPWR VDPWR VGND net126 net132 sky130_fd_sc_hd__clkbuf_4
X_2587_ VGND VDPWR VDPWR VGND net21 net174 _0101_ clknet_leaf_6_clk sky130_fd_sc_hd__dfrtp_1
Xfanout137 VDPWR VGND VDPWR VGND net138 net137 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout148 VGND VDPWR VDPWR VGND net148 _1173_ sky130_fd_sc_hd__clkbuf_4
X_1469_ VDPWR VGND VDPWR VGND net266 dig_ctrl_inst.spi_data_o\[4\] dig_ctrl_inst.data_out\[4\]
+ _0164_ _1162_ sky130_fd_sc_hd__a22o_1
Xfanout159 VGND VDPWR VDPWR VGND net159 _1152_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_3 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
X_1607_ VGND VDPWR VDPWR VGND net130 net120 net101 _0272_ sky130_fd_sc_hd__and3_4
Xfanout115 VGND VDPWR VDPWR VGND _1176_ net115 sky130_fd_sc_hd__clkbuf_2
X_1538_ VGND VDPWR VDPWR VGND _0208_ _0185_ _0206_ _0207_ sky130_fd_sc_hd__a21bo_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[45\].gen_latches\[0\].p_latch VGND VDPWR
+ VDPWR VGND net242 dig_ctrl_inst.latch_mem_inst.gclk\[45\] dig_ctrl_inst.latch_mem_inst.RAM\[45\]\[0\]
+ sky130_fd_sc_hd__dlxtp_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[0\].gen_latches\[4\].p_latch VGND VDPWR VDPWR
+ VGND net206 dig_ctrl_inst.latch_mem_inst.gclk\[0\] dig_ctrl_inst.latch_mem_inst.RAM\[0\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_0_3 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
Xdig_ctrl_inst.latch_mem_inst.gen_words\[33\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND net180 dig_ctrl_inst.latch_mem_inst.gclk\[33\] dig_ctrl_inst.latch_mem_inst.RAM\[33\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
X_2510_ VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.data\[1\] net153 _0036_ clknet_leaf_10_clk
+ sky130_fd_sc_hd__dfrtp_1
X_2441_ VGND VDPWR VDPWR VGND _0107_ dig_ctrl_inst.spi_addr\[0\] _1024_ _1025_ sky130_fd_sc_hd__o21a_1
X_1323_ VDPWR VGND VDPWR VGND net259 _1165_ net263 dig_ctrl_inst.cpu_inst.regs\[3\]\[4\]
+ sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[22\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND net199 dig_ctrl_inst.latch_mem_inst.gclk\[22\] dig_ctrl_inst.latch_mem_inst.RAM\[22\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_59_35 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2372_ VGND VDPWR VDPWR VGND _1069_ _0189_ _0769_ _1002_ sky130_fd_sc_hd__and3_4
XFILLER_0_11_249 VGND VDPWR VDPWR VGND sky130_ef_sc_hd__decap_12
Xdig_ctrl_inst.latch_mem_inst.gen_words\[11\].gen_latches\[3\].p_latch VGND VDPWR
+ VDPWR VGND net217 dig_ctrl_inst.latch_mem_inst.gclk\[11\] dig_ctrl_inst.latch_mem_inst.RAM\[11\]\[3\]
+ sky130_fd_sc_hd__dlxtp_1
X_1254_ VDPWR VGND VDPWR VGND _1094_ _1063_ _1096_ _1093_ _1095_ sky130_fd_sc_hd__or4_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[49\].gen_latches\[1\].p_latch VGND VDPWR
+ VDPWR VGND net232 dig_ctrl_inst.latch_mem_inst.gclk\[49\] dig_ctrl_inst.latch_mem_inst.RAM\[49\]\[1\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_20_29 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[4\].gen_latches\[5\].p_latch VGND VDPWR VDPWR
+ VGND net198 dig_ctrl_inst.latch_mem_inst.gclk\[4\] dig_ctrl_inst.latch_mem_inst.RAM\[4\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
X_1941_ VGND VDPWR VDPWR VGND _0601_ net90 dig_ctrl_inst.latch_mem_inst.RAM\[43\]\[5\]
+ net108 net57 sky130_fd_sc_hd__and4_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[26\].gen_latches\[6\].p_latch VGND VDPWR
+ VDPWR VGND net192 dig_ctrl_inst.latch_mem_inst.gclk\[26\] dig_ctrl_inst.latch_mem_inst.RAM\[26\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
X_1872_ VGND VDPWR VDPWR VGND _0533_ net102 dig_ctrl_inst.latch_mem_inst.RAM\[37\]\[4\]
+ net119 net54 sky130_fd_sc_hd__and4_1
X_2424_ VGND VDPWR VDPWR VGND net139 dig_ctrl_inst.cpu_inst.port_o\[6\] net328 _0102_
+ sky130_fd_sc_hd__mux2_1
X_1306_ VGND VDPWR VDPWR VGND net263 net259 _1148_ dig_ctrl_inst.cpu_inst.regs\[2\]\[5\]
+ sky130_fd_sc_hd__and3b_1
X_2286_ VGND VDPWR VDPWR VGND _0927_ _0767_ _0926_ _0928_ _0768_ sky130_fd_sc_hd__a2bb2o_1
X_2355_ VGND VDPWR VDPWR VGND _0991_ _0992_ net352 _0054_ sky130_fd_sc_hd__mux2_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[15\].gen_latches\[4\].p_latch VGND VDPWR
+ VDPWR VGND net203 dig_ctrl_inst.latch_mem_inst.gclk\[15\] dig_ctrl_inst.latch_mem_inst.RAM\[15\]\[4\]
+ sky130_fd_sc_hd__dlxtp_1
X_1237_ VGND VDPWR VDPWR VGND _1079_ _1038_ _1063_ dig_ctrl_inst.cpu_inst.regs\[1\]\[0\]
+ _1077_ sky130_fd_sc_hd__a211o_1
XFILLER_0_19_113 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.genblk1\[29\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[29\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[29\]._gclk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_193 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
Xdig_ctrl_inst.latch_mem_inst.gen_words\[8\].gen_latches\[6\].p_latch VGND VDPWR VDPWR
+ VGND net191 dig_ctrl_inst.latch_mem_inst.gclk\[8\] dig_ctrl_inst.latch_mem_inst.RAM\[8\]\[6\]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_0_249 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
X_2140_ VGND VDPWR VDPWR VGND _0785_ net149 _0784_ _0786_ sky130_fd_sc_hd__o21ai_1
X_2071_ VGND VDPWR VDPWR VGND _0729_ net106 dig_ctrl_inst.latch_mem_inst.RAM\[11\]\[7\]
+ net127 net91 sky130_fd_sc_hd__and4_1
X_1924_ VDPWR VGND VDPWR VGND net129 _0584_ dig_ctrl_inst.latch_mem_inst.RAM\[6\]\[5\]
+ net95 sky130_fd_sc_hd__and3_2
X_1855_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[2\]\[3\] _1178_ _0517_
+ dig_ctrl_inst.latch_mem_inst.RAM\[25\]\[3\] _0129_ sky130_fd_sc_hd__a22o_1
X_1786_ VGND VDPWR VDPWR VGND _0449_ net121 dig_ctrl_inst.latch_mem_inst.RAM\[17\]\[2\]
+ net137 net68 sky130_fd_sc_hd__and4_1
Xdig_ctrl_inst.latch_mem_inst.gen_words\[19\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND net196 dig_ctrl_inst.latch_mem_inst.gclk\[19\] dig_ctrl_inst.latch_mem_inst.RAM\[19\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
X_2407_ VGND VDPWR VDPWR VGND _0176_ net350 dig_ctrl_inst.spi_data_o\[6\] _0087_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_3 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_6
X_2338_ VGND VDPWR VDPWR VGND _0172_ _0808_ _0806_ _0977_ sky130_fd_sc_hd__mux2_1
X_2269_ VGND VDPWR VDPWR VGND _0858_ _0911_ _0910_ _0787_ _0857_ _0795_ sky130_fd_sc_hd__o221ai_1
Xhold40 VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_data_i\[1\] net322 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_141 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_8
Xhold51 VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[2\]\[7\] net333 sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[1\]\[7\] net344 sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 VGND VDPWR VDPWR VGND dig_ctrl_inst.cpu_inst.regs\[0\]\[7\] net355 sky130_fd_sc_hd__dlygate4sd3_1
Xdig_ctrl_inst.latch_mem_inst.genblk1\[11\].clock_gate VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.data_we\[11\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[11\]._gclk clknet_leaf_18_clk sky130_fd_sc_hd__dlclkp_1
XANTENNA_4 VGND VDPWR VDPWR VGND _0325_ sky130_fd_sc_hd__diode_2
XFILLER_0_67_57 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
X_1640_ VDPWR VGND VDPWR VGND _0299_ _0305_ _0300_ _0304_ sky130_fd_sc_hd__or3_1
X_1571_ VGND VDPWR VDPWR VGND _0237_ net163 _1114_ sky130_fd_sc_hd__nand2_1
X_2123_ VGND VDPWR VDPWR VGND _0769_ _0766_ _0767_ sky130_fd_sc_hd__nand2b_1
X_2054_ VGND VDPWR VDPWR VGND _0712_ net89 dig_ctrl_inst.latch_mem_inst.RAM\[27\]\[7\]
+ net104 net59 sky130_fd_sc_hd__and4_1
X_1838_ VDPWR VGND VDPWR VGND dig_ctrl_inst.latch_mem_inst.RAM\[37\]\[3\] _0140_ _0500_
+ dig_ctrl_inst.latch_mem_inst.RAM\[53\]\[3\] _0154_ sky130_fd_sc_hd__a22o_1
X_1907_ VGND VDPWR VDPWR VGND _0529_ _0568_ _0536_ dig_ctrl_inst.latch_mem_inst.RAM\[23\]\[4\]
+ _0128_ _0534_ sky130_fd_sc_hd__a2111o_1
X_1769_ VGND VDPWR VDPWR VGND _0429_ _0432_ _0431_ dig_ctrl_inst.latch_mem_inst.RAM\[7\]\[2\]
+ _1184_ _0430_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_12_141 VDPWR VGND VDPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_35_233 VGND VDPWR VDPWR VGND sky130_fd_sc_hd__decap_4
Xoutput30 VDPWR VGND VDPWR VGND uo_out[5] net30 sky130_fd_sc_hd__buf_2
Xdig_ctrl_inst.latch_mem_inst.genblk1\[9\].clock_buffer VGND VDPWR VDPWR VGND dig_ctrl_inst.latch_mem_inst.gclk\[9\]
+ dig_ctrl_inst.latch_mem_inst.genblk1\[9\]._gclk sky130_fd_sc_hd__clkbuf_4
Xdig_ctrl_inst.latch_mem_inst.gen_words\[63\].gen_latches\[7\].p_latch VGND VDPWR
+ VDPWR VGND net184 dig_ctrl_inst.latch_mem_inst.gclk\[63\] dig_ctrl_inst.latch_mem_inst.RAM\[63\]\[7\]
+ sky130_fd_sc_hd__dlxtp_1
X_1485_ VGND VDPWR VDPWR VGND dig_ctrl_inst.spi_receiver_inst.spi_cs_sync dig_ctrl_inst.spi_receiver_inst.spi_sclk_sync
+ dig_ctrl_inst.spi_receiver_inst.spi_sclk_delayed _0176_ sky130_fd_sc_hd__or3b_4
X_1554_ VDPWR VGND VDPWR VGND _0220_ dig_ctrl_inst.cpu_inst.regs\[1\]\[7\] _1035_
+ _1068_ dig_ctrl_inst.cpu_inst.regs\[2\]\[7\] net177 sky130_fd_sc_hd__a221o_1
X_1623_ VDPWR VGND VDPWR VGND net86 _0288_ dig_ctrl_inst.latch_mem_inst.RAM\[24\]\[0\]
+ net66 sky130_fd_sc_hd__and3_2
Xdig_ctrl_inst.latch_mem_inst.gen_words\[52\].gen_latches\[5\].p_latch VGND VDPWR
+ VDPWR VGND net197 dig_ctrl_inst.latch_mem_inst.gclk\[52\] dig_ctrl_inst.latch_mem_inst.RAM\[52\]\[5\]
+ sky130_fd_sc_hd__dlxtp_1
.ends

.subckt res_poly a_n141_4996# a_n141_n5432# VSUBS
X0 a_n141_4996# a_n141_n5432# VSUBS sky130_fd_pr__res_high_po_1p41 l=50.12
.ends

.subckt sky130_leo_ip__rdac_8bit D0 D1 D2 D3 D4 D5 D6 D7 OUT VGND
Xres_poly_0 m1_5556_10930# m1_4470_10930# VGND res_poly
Xres_poly_1 m1_4470_10930# m1_4832_499# VGND res_poly
Xres_poly_2 m1_4470_10930# m1_3384_10930# VGND res_poly
Xres_poly_3 D2 m1_3746_499# VGND res_poly
Xres_poly_4 m1_3384_10930# m1_3746_499# VGND res_poly
Xres_poly_5 m1_3384_10930# m1_2298_10930# VGND res_poly
Xres_poly_6 D1 m1_2660_499# VGND res_poly
Xres_poly_7 m1_2298_10930# m1_2660_499# VGND res_poly
Xres_poly_8 m1_2298_10930# m1_1212_10930# VGND res_poly
Xres_poly_9 VGND m1_1574_499# VGND res_poly
Xres_poly_21 D6 m1_8090_499# VGND res_poly
Xres_poly_20 m1_7728_10930# m1_8090_499# VGND res_poly
Xres_poly_10 m1_1212_10930# m1_1574_499# VGND res_poly
Xres_poly_22 OUT m1_7728_10930# VGND res_poly
Xres_poly_11 m1_1212_10930# m1_850_499# VGND res_poly
Xres_poly_23 OUT m1_9176_499# VGND res_poly
Xres_poly_12 VGND VGND VGND res_poly
Xres_poly_24 D7 m1_9176_499# VGND res_poly
Xres_poly_13 D3 m1_4832_499# VGND res_poly
Xres_poly_25 VGND VGND VGND res_poly
Xres_poly_14 m1_5556_10930# m1_5918_499# VGND res_poly
Xres_poly_15 D4 m1_5918_499# VGND res_poly
Xres_poly_26 D0 m1_850_499# VGND res_poly
Xres_poly_16 m1_6642_10930# m1_5556_10930# VGND res_poly
Xres_poly_18 D5 m1_7004_499# VGND res_poly
Xres_poly_17 m1_6642_10930# m1_7004_499# VGND res_poly
Xres_poly_19 m1_7728_10930# m1_6642_10930# VGND res_poly
.ends

.subckt pfet a_60_n40# w_n242_n247# a_160_0# a_0_0#
X0 a_160_0# a_60_n40# a_0_0# w_n242_n247# sky130_fd_pr__pfet_g5v0d10v5 ad=6 pd=40.6 as=6 ps=40.6 w=20 l=0.5
.ends

.subckt res_poly$1 a_n285_2496# a_n415_n3062# a_n285_n2932#
X0 a_n285_2496# a_n285_n2932# a_n415_n3062# sky130_fd_pr__res_xhigh_po_2p85 l=25.12
.ends

.subckt pfet$10 a_60_n40# w_n242_n247# a_1060_0# a_0_0#
X0 a_1060_0# a_60_n40# a_0_0# w_n242_n247# sky130_fd_pr__pfet_g5v0d10v5 ad=3 pd=20.6 as=3 ps=20.6 w=10 l=5
.ends

.subckt nfet$5 a_60_n40# a_160_0# a_0_0# a_n149_n154#
X0 a_160_0# a_60_n40# a_0_0# a_n149_n154# sky130_fd_pr__nfet_g5v0d10v5 ad=0.3 pd=2.6 as=0.3 ps=2.6 w=1 l=0.5
.ends

.subckt pfet$9 a_60_n40# w_n242_n247# a_1060_0# a_0_0#
X0 a_1060_0# a_60_n40# a_0_0# w_n242_n247# sky130_fd_pr__pfet_g5v0d10v5 ad=0.3 pd=2.6 as=0.3 ps=2.6 w=1 l=5
.ends

.subckt sky130_fd_sc_hvl__buf_4$VAR1 VPB VPWR VNB VGND A X
X0 a_149_81# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.21 ps=1.78 w=1.5 l=0.5
X1 VGND a_149_81# X VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X2 X a_149_81# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.21375 ps=2.07 w=0.75 l=0.5
X3 X a_149_81# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X4 VPWR a_149_81# X VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X5 a_149_81# A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.105 ps=1.03 w=0.75 l=0.5
X6 VPWR a_149_81# X VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X7 X a_149_81# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.4275 ps=3.57 w=1.5 l=0.5
X8 X a_149_81# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X9 VGND a_149_81# X VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
.ends

.subckt pfet$5 a_60_n40# w_n242_n247# a_160_0# a_0_0#
X0 a_160_0# a_60_n40# a_0_0# w_n242_n247# sky130_fd_pr__pfet_g5v0d10v5 ad=1.5 pd=10.6 as=1.5 ps=10.6 w=5 l=0.5
.ends

.subckt sky130_fd_sc_hvl__buf_4$1 VPB VPWR VNB VGND A X
X0 a_149_81# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.21 ps=1.78 w=1.5 l=0.5
X1 VGND a_149_81# X VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X2 X a_149_81# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.21375 ps=2.07 w=0.75 l=0.5
X3 X a_149_81# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X4 VPWR a_149_81# X VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X5 a_149_81# A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.105 ps=1.03 w=0.75 l=0.5
X6 VPWR a_149_81# X VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X7 X a_149_81# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.4275 ps=3.57 w=1.5 l=0.5
X8 X a_149_81# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X9 VGND a_149_81# X VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
.ends

.subckt nfet$6 a_60_n40# a_160_0# a_0_0# a_n149_n154#
X0 a_160_0# a_60_n40# a_0_0# a_n149_n154# sky130_fd_pr__nfet_g5v0d10v5 ad=3 pd=20.6 as=3 ps=20.6 w=10 l=0.5
.ends

.subckt nfet$4 a_60_n40# a_160_0# a_0_0# a_n149_n154#
X0 a_160_0# a_60_n40# a_0_0# a_n149_n154# sky130_fd_pr__nfet_g5v0d10v5 ad=1.5 pd=10.6 as=1.5 ps=10.6 w=5 l=0.5
.ends

.subckt sky130_fd_sc_hvl__nand2_1 VPB VPWR VNB VGND B Y A
X0 a_233_111# B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.07875 pd=0.96 as=0.21375 ps=2.07 w=0.75 l=0.5
X1 Y A a_233_111# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.07875 ps=0.96 w=0.75 l=0.5
X2 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.21 ps=1.78 w=1.5 l=0.5
X3 Y B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.4275 ps=3.57 w=1.5 l=0.5
.ends

.subckt sky130_leo_ip__comparator VDD IN_P OUT_P IN_N CLK_N OUT_N VSS
Xpfet_0 IN_N VDD m1_1831_3328# COMP_N pfet
Xpfet_1 IN_P VDD COMP_P m1_1831_3328# pfet
Xres_poly$1_0 m1_282_7668# VSS VSS res_poly$1
Xpfet$10_0 m1_282_7668# VDD VDD m1_1831_3328# pfet$10
Xnfet$5_0 COMP_P SR_reset VSS VSS nfet$5
Xnfet$5_1 COMP_N SR_set VSS VSS nfet$5
Xpfet$9_0 m1_282_7668# VDD m1_282_7668# VDD pfet$9
Xsky130_fd_sc_hvl__buf_4$VAR1_0 VDD VDD VSS VSS sky130_fd_sc_hvl__nand2_1_1/Y OUT_N
+ sky130_fd_sc_hvl__buf_4$VAR1
Xpfet$5_0 COMP_P VDD VDD SR_reset pfet$5
Xsky130_fd_sc_hvl__buf_4$1_0 VDD VDD VSS VSS sky130_fd_sc_hvl__nand2_1_1/A OUT_P sky130_fd_sc_hvl__buf_4$1
Xpfet$5_1 COMP_N VDD VDD SR_set pfet$5
Xnfet$6_0 CLK_N COMP_P COMP_N VSS nfet$6
Xnfet$4_0 COMP_N VSS COMP_P VSS nfet$4
Xsky130_fd_sc_hvl__nand2_1_0 VDD VDD VSS VSS sky130_fd_sc_hvl__nand2_1_1/Y sky130_fd_sc_hvl__nand2_1_1/A
+ SR_reset sky130_fd_sc_hvl__nand2_1
Xnfet$4_1 COMP_P COMP_N VSS VSS nfet$4
Xsky130_fd_sc_hvl__nand2_1_1 VDD VDD VSS VSS SR_set sky130_fd_sc_hvl__nand2_1_1/Y
+ sky130_fd_sc_hvl__nand2_1_1/A sky130_fd_sc_hvl__nand2_1
.ends

.subckt tt_um_tt08_aicd_playground VAPWR ui_in[7] ui_in[6] ui_in[5] ui_in[4] ui_in[3]
+ ui_in[2] ui_in[1] ui_in[0] VDPWR VGND uio_in[7] uio_in[6] uio_in[5] uio_in[4] uio_in[3]
+ uio_in[2] uio_in[1] uio_in[0] ena uo_out[7] uo_out[6] uo_out[5] uo_out[4] uo_out[3]
+ uo_out[2] uo_out[1] uo_out[0] clk rst_n uio_out[7] uio_out[6] uio_out[5] uio_out[4]
+ uio_out[3] uio_out[2] uio_out[1] uio_out[0] uio_oe[7] uio_oe[6] uio_oe[5] uio_oe[4]
+ uio_oe[3] uio_oe[2] uio_oe[1] uio_oe[0] ua[7] ua[6] ua[5] ua[4] ua[3] ua[2] ua[1]
+ ua[0]
Xsky130_leo_ip__levelshifter_up_1 VAPWR VDPWR sky130_fd_sc_hvl__buf_4_1/A dig_ctrl_top_0/port_ms_o[6]
+ VGND sky130_leo_ip__levelshifter_up
Xsky130_leo_ip__levelshifter_up_2 VAPWR VDPWR sky130_fd_sc_hvl__buf_4_2/A dig_ctrl_top_0/port_ms_o[5]
+ VGND sky130_leo_ip__levelshifter_up
Xsky130_leo_ip__levelshifter_up_3 VAPWR VDPWR sky130_fd_sc_hvl__buf_4_3/A dig_ctrl_top_0/port_ms_o[4]
+ VGND sky130_leo_ip__levelshifter_up
Xsky130_leo_ip__levelshifter_up_4 VAPWR VDPWR sky130_fd_sc_hvl__buf_4_4/A dig_ctrl_top_0/port_ms_o[3]
+ VGND sky130_leo_ip__levelshifter_up
Xsky130_leo_ip__levelshifter_up_5 VAPWR VDPWR sky130_fd_sc_hvl__buf_4_5/A dig_ctrl_top_0/port_ms_o[2]
+ VGND sky130_leo_ip__levelshifter_up
Xsky130_leo_ip__levelshifter_up_6 VAPWR VDPWR sky130_fd_sc_hvl__buf_4_6/A dig_ctrl_top_0/port_ms_o[1]
+ VGND sky130_leo_ip__levelshifter_up
Xsky130_fd_sc_hvl__buf_4_0 VGND VGND VAPWR VAPWR sky130_fd_sc_hvl__buf_4_0/X sky130_fd_sc_hvl__buf_4_0/A
+ sky130_fd_sc_hvl__buf_4
Xsky130_leo_ip__levelshifter_up_7 VAPWR VDPWR sky130_fd_sc_hvl__buf_4_7/A dig_ctrl_top_0/port_ms_o[0]
+ VGND sky130_leo_ip__levelshifter_up
Xsky130_fd_sc_hvl__buf_4_1 VGND VGND VAPWR VAPWR sky130_fd_sc_hvl__buf_4_1/X sky130_fd_sc_hvl__buf_4_1/A
+ sky130_fd_sc_hvl__buf_4
Xsky130_fd_sc_hvl__buf_4_2 VGND VGND VAPWR VAPWR sky130_fd_sc_hvl__buf_4_2/X sky130_fd_sc_hvl__buf_4_2/A
+ sky130_fd_sc_hvl__buf_4
Xsky130_leo_ip__levelshifter_down_0 dig_ctrl_top_0/port_ms_i sky130_leo_ip__comparator_0/OUT_P
+ VGND VDPWR sky130_leo_ip__levelshifter_down
Xdig_ctrl_top_0 clk ena rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5]
+ uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7]
+ uio_oe[0] uio_oe[1] uio_oe[3] uio_oe[4] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1]
+ uio_out[2] uio_out[3] uio_out[4] uio_out[6] uio_out[7] uo_out[0] uo_out[1] uo_out[2]
+ uo_out[3] uo_out[4] uo_out[5] uo_out[6] uo_out[7] dig_ctrl_top_0/clk_o dig_ctrl_top_0/port_ms_i
+ dig_ctrl_top_0/port_ms_o[0] dig_ctrl_top_0/port_ms_o[1] dig_ctrl_top_0/port_ms_o[2]
+ dig_ctrl_top_0/port_ms_o[3] dig_ctrl_top_0/port_ms_o[4] dig_ctrl_top_0/port_ms_o[5]
+ dig_ctrl_top_0/port_ms_o[6] dig_ctrl_top_0/port_ms_o[7] uio_out[5] ui_in[6] uio_oe[5]
+ uio_oe[2] ui_in[7] VGND VDPWR dig_ctrl_top
Xsky130_fd_sc_hvl__buf_4_3 VGND VGND VAPWR VAPWR sky130_fd_sc_hvl__buf_4_3/X sky130_fd_sc_hvl__buf_4_3/A
+ sky130_fd_sc_hvl__buf_4
Xsky130_fd_sc_hvl__buf_4_4 VGND VGND VAPWR VAPWR sky130_fd_sc_hvl__buf_4_4/X sky130_fd_sc_hvl__buf_4_4/A
+ sky130_fd_sc_hvl__buf_4
Xsky130_fd_sc_hvl__buf_4_5 VGND VGND VAPWR VAPWR sky130_fd_sc_hvl__buf_4_5/X sky130_fd_sc_hvl__buf_4_5/A
+ sky130_fd_sc_hvl__buf_4
Xsky130_fd_sc_hvl__buf_4_6 VGND VGND VAPWR VAPWR sky130_fd_sc_hvl__buf_4_6/X sky130_fd_sc_hvl__buf_4_6/A
+ sky130_fd_sc_hvl__buf_4
Xsky130_fd_sc_hvl__buf_4_7 VGND VGND VAPWR VAPWR sky130_fd_sc_hvl__buf_4_7/X sky130_fd_sc_hvl__buf_4_7/A
+ sky130_fd_sc_hvl__buf_4
Xsky130_leo_ip__rdac_8bit_0 sky130_fd_sc_hvl__buf_4_7/X sky130_fd_sc_hvl__buf_4_6/X
+ sky130_fd_sc_hvl__buf_4_5/X sky130_fd_sc_hvl__buf_4_4/X sky130_fd_sc_hvl__buf_4_3/X
+ sky130_fd_sc_hvl__buf_4_2/X sky130_fd_sc_hvl__buf_4_1/X sky130_fd_sc_hvl__buf_4_0/X
+ ua[1] VGND sky130_leo_ip__rdac_8bit
Xsky130_leo_ip__comparator_0 VAPWR ua[0] sky130_leo_ip__comparator_0/OUT_P ua[1] dig_ctrl_top_0/clk_o
+ sky130_leo_ip__comparator_0/OUT_N VGND sky130_leo_ip__comparator
Xsky130_leo_ip__levelshifter_up_0 VAPWR VDPWR sky130_fd_sc_hvl__buf_4_0/A dig_ctrl_top_0/port_ms_o[7]
+ VGND sky130_leo_ip__levelshifter_up
.ends

